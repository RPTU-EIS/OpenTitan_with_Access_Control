function automatic clk_gating_disabled();
    clk_gating_disabled = (
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.clock_en &&
        top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.clock_en
    );
endfunction

function automatic input_equivalence_rv_core_ibex();
    input_equivalence_rv_core_ibex = (
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.clk_i              == top_level_upec.top_earlgrey_1.u_rv_core_ibex.clk_i               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.rst_ni             == top_level_upec.top_earlgrey_1.u_rv_core_ibex.rst_ni              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.clk_esc_i          == top_level_upec.top_earlgrey_1.u_rv_core_ibex.clk_esc_i       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.rst_esc_ni         == top_level_upec.top_earlgrey_1.u_rv_core_ibex.rst_esc_ni      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.ram_cfg_i          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.ram_cfg_i       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.hart_id_i          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.hart_id_i       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.boot_addr_i        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.boot_addr_i     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_i_i             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_i_i          &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_d_i             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_d_i          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.irq_software_i     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.irq_software_i  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.irq_timer_i        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.irq_timer_i     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.irq_external_i     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.irq_external_i  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.esc_tx_i           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.esc_tx_i        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.debug_req_i        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.debug_req_i     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.lc_cpu_en_i        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.lc_cpu_en_i     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.pwrmgr_cpu_en_i    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.pwrmgr_cpu_en_i &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.scan_rst_ni        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.scan_rst_ni     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.scanmode_i         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.scanmode_i
    );
endfunction

function automatic output_equivalence_rv_core_ibex();
    output_equivalence_rv_core_ibex = (
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_i_o         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_i_o          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_d_o         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_d_o          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.esc_rx_o       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.esc_rx_o        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.crash_dump_o   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.crash_dump_o    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.core_sleep_o   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.core_sleep_o
    );
endfunction

function automatic visible_soc_state_equivalence_rv_core_ibex();
    visible_soc_state_equivalence_rv_core_ibex = (
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstatus_csr.rdata_q                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstatus_csr.rdata_q                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mie_csr.rdata_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mie_csr.rdata_q                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtvec_csr.rdata_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtvec_csr.rdata_q                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcountinhibit_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcountinhibit_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mscratch_csr.rdata_q                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mscratch_csr.rdata_q                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mepc_csr.rdata_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mepc_csr.rdata_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mcause_csr.rdata_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mcause_csr.rdata_q                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtval_csr.rdata_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtval_csr.rdata_q                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.irq_software_i                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.irq_software_i                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.irq_timer_i                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.irq_timer_i                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.irq_external_i                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.irq_external_i                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.irq_fast_i                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.irq_fast_i                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_cfg_csr.rdata_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_cfg_csr.rdata_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_cfg_csr.rdata_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_cfg_csr.rdata_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_cfg_csr.rdata_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_cfg_csr.rdata_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_cfg_csr.rdata_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_cfg_csr.rdata_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_cfg_csr.rdata_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_cfg_csr.rdata_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_cfg_csr.rdata_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_cfg_csr.rdata_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_cfg_csr.rdata_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_cfg_csr.rdata_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_cfg_csr.rdata_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_cfg_csr.rdata_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_cfg_csr.rdata_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_cfg_csr.rdata_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_cfg_csr.rdata_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_cfg_csr.rdata_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_cfg_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_cfg_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_cfg_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_cfg_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_cfg_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_cfg_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_cfg_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_cfg_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_cfg_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_cfg_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_cfg_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_cfg_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_addr_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_addr_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_addr_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_addr_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_addr_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_addr_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_addr_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_addr_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_addr_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_addr_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_addr_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_addr_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_addr_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_addr_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_addr_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_addr_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_addr_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_addr_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_addr_csr.rdata_q     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_addr_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_addr_csr.rdata_q    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_addr_csr.rdata_q &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_addr_csr.rdata_q    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_addr_csr.rdata_q &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_addr_csr.rdata_q    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_addr_csr.rdata_q &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_addr_csr.rdata_q    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_addr_csr.rdata_q &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_addr_csr.rdata_q    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_addr_csr.rdata_q &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_addr_csr.rdata_q    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_addr_csr.rdata_q &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.u_pmp_mseccfg.rdata_q                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.u_pmp_mseccfg.rdata_q                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.u_tselect_csr.rdata_q                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.u_tselect_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.selected_tmatch_control                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.selected_tmatch_control              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.selected_tmatch_value                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.selected_tmatch_value                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dcsr_csr.rdata_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dcsr_csr.rdata_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_depc_csr.rdata_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_depc_csr.rdata_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch0_csr.rdata_q                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch0_csr.rdata_q                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch1_csr.rdata_q                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch1_csr.rdata_q                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_cpuctrl_csr.rdata_q                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_cpuctrl_csr.rdata_q                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcycle_counter_i.counter_q                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcycle_counter_i.counter_q                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.minstret_counter_i.counter_q                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.minstret_counter_i.counter_q                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[0].gen_imp.mcounters_variable_i.counter_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[0].gen_imp.mcounters_variable_i.counter_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[1].gen_imp.mcounters_variable_i.counter_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[1].gen_imp.mcounters_variable_i.counter_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[2].gen_imp.mcounters_variable_i.counter_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[2].gen_imp.mcounters_variable_i.counter_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[3].gen_imp.mcounters_variable_i.counter_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[3].gen_imp.mcounters_variable_i.counter_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[4].gen_imp.mcounters_variable_i.counter_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[4].gen_imp.mcounters_variable_i.counter_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[5].gen_imp.mcounters_variable_i.counter_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[5].gen_imp.mcounters_variable_i.counter_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[6].gen_imp.mcounters_variable_i.counter_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[6].gen_imp.mcounters_variable_i.counter_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[7].gen_imp.mcounters_variable_i.counter_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[7].gen_imp.mcounters_variable_i.counter_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[8].gen_imp.mcounters_variable_i.counter_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[8].gen_imp.mcounters_variable_i.counter_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[9].gen_imp.mcounters_variable_i.counter_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[9].gen_imp.mcounters_variable_i.counter_q   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_regfile_ff.register_file_i.rf_reg_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_regfile_ff.register_file_i.rf_reg_q
        );
endfunction

function automatic micro_soc_state_equivalence_rv_core_ibex();
    micro_soc_state_equivalence_rv_core_ibex = (
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_d_ibex.g_multiple_reqs.source_q                                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_d_ibex.g_multiple_reqs.source_q                                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_d_ibex.intg_err_q                                                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_d_ibex.intg_err_q                                                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_d_ibex.outstanding_reqs_q                                                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_d_ibex.outstanding_reqs_q                                                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_i_ibex.g_multiple_reqs.source_q                                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_i_ibex.g_multiple_reqs.source_q                                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_i_ibex.intg_err_q                                                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_i_ibex.intg_err_q                                                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_i_ibex.outstanding_reqs_q                                                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_i_ibex.outstanding_reqs_q                                                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.core_busy_q                                                                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.core_busy_q                                                                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.core_clock_gate_i.gen_generic.u_impl_generic.en_latch                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.core_clock_gate_i.gen_generic.u_impl_generic.en_latch                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.fetch_enable_q                                                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.fetch_enable_q                                                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.core_outputs_q                                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.core_outputs_q                                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.rst_shadow_cnt_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.rst_shadow_cnt_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.rst_shadow_set_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.rst_shadow_set_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_data_rdata_q                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_data_rdata_q                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_inputs_q                                                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_inputs_q                                                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_tag_rdata_q                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_tag_rdata_q                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.u_pmp_mseccfg.rdata_q                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.u_pmp_mseccfg.rdata_q                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[0].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[0].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[1].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[1].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[2].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[2].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[3].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[3].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[4].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[4].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[5].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[5].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[6].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[6].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[7].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[7].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[8].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[8].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[9].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[9].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr.rdata_q == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr.rdata_q   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr.rdata_q    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.u_tselect_csr.rdata_q                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.u_tselect_csr.rdata_q                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.mcountinhibit_q                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.mcountinhibit_q                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.mcycle_counter_i.counter_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.mcycle_counter_i.counter_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.minstret_counter_i.counter_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.minstret_counter_i.counter_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.priv_lvl_q                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.priv_lvl_q                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_cpuctrl_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_cpuctrl_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dcsr_csr.rdata_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dcsr_csr.rdata_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_depc_csr.rdata_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_depc_csr.rdata_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dscratch0_csr.rdata_q                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dscratch0_csr.rdata_q                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dscratch1_csr.rdata_q                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dscratch1_csr.rdata_q                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mcause_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mcause_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mepc_csr.rdata_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mepc_csr.rdata_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mie_csr.rdata_q                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mie_csr.rdata_q                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mscratch_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mscratch_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_cause_csr.rdata_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_cause_csr.rdata_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_epc_csr.rdata_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_epc_csr.rdata_q                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstatus_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstatus_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mtval_csr.rdata_q                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mtval_csr.rdata_q                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mtvec_csr.rdata_q                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mtvec_csr.rdata_q                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_single_cycle.mult_state_q         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_single_cycle.mult_state_q          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.branch_jump_set_done_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.branch_jump_set_done_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.ctrl_fsm_cs                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.ctrl_fsm_cs                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.debug_mode_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.debug_mode_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.do_single_step_q                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.do_single_step_q                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.enter_debug_mode_prio_q                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.enter_debug_mode_prio_q                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exc_req_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exc_req_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exception_req_accepted                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exception_req_accepted                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exception_req_pending                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exception_req_pending                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.expect_exception_pc_set                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.expect_exception_pc_set                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.illegal_insn_q                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.illegal_insn_q                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.load_err_q                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.load_err_q                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.nmi_mode_q                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.nmi_mode_q                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.seen_exception_pc_set                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.seen_exception_pc_set                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.store_err_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.store_err_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.g_branch_set_flop.branch_set_raw_q                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.g_branch_set_flop.branch_set_raw_q                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.g_sec_branch_taken.branch_taken_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.g_sec_branch_taken.branch_taken_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.id_fsm_q                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.id_fsm_q                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.imd_val_q                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.imd_val_q                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.dummy_instr_id_o                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.dummy_instr_id_o                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.g_secure_pc.prev_instr_seq_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.g_secure_pc.prev_instr_seq_q                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_cnt_q                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_cnt_q                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_instr_seed_q                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_instr_seed_q                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.cnt_q            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.cnt_q             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.perturbed_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.perturbed_q       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.lfsr_q                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.lfsr_q                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_addr_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_addr_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_busy_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_busy_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_cache_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_cache_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_data_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_data_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_err_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_err_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_cnt_q                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_cnt_q                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_done_q                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_done_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_hold_q                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_hold_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_hit_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_hit_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_in_ic1                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_in_ic1                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_older_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_older_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_out_cnt_q                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_out_cnt_q                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ram_done_q                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ram_done_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_rvd_cnt_q                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_rvd_cnt_q                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_stale_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_stale_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_way_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_way_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_index_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_index_q       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_ways_q       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_ways_q        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_write_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_write_q       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.lookup_index_ic1            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.lookup_index_ic1             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.inval_index_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.inval_index_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.inval_prog_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.inval_prog_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.lookup_addr_ic1                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.lookup_addr_ic1                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.lookup_valid_ic1                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.lookup_valid_ic1                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.output_addr_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.output_addr_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.prefetch_addr_q                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.prefetch_addr_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.reset_inval_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.reset_inval_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.round_robin_way_q                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.round_robin_way_q                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_data_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_data_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_err_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_err_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_valid_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_valid_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.illegal_c_insn_id_o                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.illegal_c_insn_id_o                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_fetch_err_o                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_fetch_err_o                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_fetch_err_plus2_o                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_fetch_err_plus2_o                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_is_compressed_id_o                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_is_compressed_id_o                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_new_id_q                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_new_id_q                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_alu_id_o                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_alu_id_o                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_c_id_o                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_c_id_o                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_id_o                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_id_o                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_valid_id_q                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_valid_id_q                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.pc_id_o                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.pc_id_o                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.addr_last_q                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.addr_last_q                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_sign_ext_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_sign_ext_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_type_q                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_type_q                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_we_q                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_we_q                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.handle_misaligned_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.handle_misaligned_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.ls_fsm_cs                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.ls_fsm_cs                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.lsu_err_q                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.lsu_err_q                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.pmp_err_q                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.pmp_err_q                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.rdata_offset_q                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.rdata_offset_q                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.rdata_q                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.rdata_q                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_waddr_wb_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_waddr_wb_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_wdata_wb_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_wdata_wb_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_we_wb_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_we_wb_q                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_compressed_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_compressed_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_count_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_count_q                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_instr_type_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_instr_type_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_pc_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_pc_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_valid_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_valid_q                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].data_bank.gen_generic.u_impl_generic.mem                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].data_bank.gen_generic.u_impl_generic.mem                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].data_bank.gen_generic.u_impl_generic.rdata_o                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].data_bank.gen_generic.u_impl_generic.rdata_o                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].tag_bank.gen_generic.u_impl_generic.mem                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].tag_bank.gen_generic.u_impl_generic.mem                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].tag_bank.gen_generic.u_impl_generic.rdata_o                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].tag_bank.gen_generic.u_impl_generic.rdata_o                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].data_bank.gen_generic.u_impl_generic.mem                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].data_bank.gen_generic.u_impl_generic.mem                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].data_bank.gen_generic.u_impl_generic.rdata_o                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].data_bank.gen_generic.u_impl_generic.rdata_o                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].tag_bank.gen_generic.u_impl_generic.mem                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].tag_bank.gen_generic.u_impl_generic.mem                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].tag_bank.gen_generic.u_impl_generic.rdata_o                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].tag_bank.gen_generic.u_impl_generic.rdata_o                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_regfile_ff.register_file_i.g_dummy_r0.rf_r0_q                                                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_regfile_ff.register_file_i.g_dummy_r0.rf_r0_q                                                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_regfile_ff.register_file_i.rf_reg_q                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_regfile_ff.register_file_i.rf_reg_q                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.u_pmp_mseccfg.rdata_q                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.u_pmp_mseccfg.rdata_q                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[0].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[0].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[1].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[1].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[2].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[2].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[3].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[3].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[4].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[4].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[5].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[5].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[6].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[6].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[7].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[7].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[8].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[8].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[9].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[9].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr.rdata_q                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr.rdata_q                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr.rdata_q                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr.rdata_q                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.u_tselect_csr.rdata_q                                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.u_tselect_csr.rdata_q                                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcountinhibit_q                                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcountinhibit_q                                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcycle_counter_i.counter_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcycle_counter_i.counter_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.minstret_counter_i.counter_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.minstret_counter_i.counter_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.priv_lvl_q                                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.priv_lvl_q                                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_cpuctrl_csr.rdata_q                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_cpuctrl_csr.rdata_q                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dcsr_csr.rdata_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dcsr_csr.rdata_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_depc_csr.rdata_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_depc_csr.rdata_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch0_csr.rdata_q                                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch0_csr.rdata_q                                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch1_csr.rdata_q                                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch1_csr.rdata_q                                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mcause_csr.rdata_q                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mcause_csr.rdata_q                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mepc_csr.rdata_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mepc_csr.rdata_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mie_csr.rdata_q                                                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mie_csr.rdata_q                                                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mscratch_csr.rdata_q                                                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mscratch_csr.rdata_q                                                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_cause_csr.rdata_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_cause_csr.rdata_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_csr.rdata_q                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_csr.rdata_q                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_epc_csr.rdata_q                                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_epc_csr.rdata_q                                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstatus_csr.rdata_q                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstatus_csr.rdata_q                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtval_csr.rdata_q                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtval_csr.rdata_q                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtvec_csr.rdata_q                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtvec_csr.rdata_q                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_single_cycle.mult_state_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_single_cycle.mult_state_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q                                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q                                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.branch_jump_set_done_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.branch_jump_set_done_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.ctrl_fsm_cs                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.ctrl_fsm_cs                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.debug_mode_q                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.debug_mode_q                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.do_single_step_q                                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.do_single_step_q                                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.enter_debug_mode_prio_q                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.enter_debug_mode_prio_q                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exc_req_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exc_req_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exception_req_accepted                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exception_req_accepted                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exception_req_pending                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exception_req_pending                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.expect_exception_pc_set                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.expect_exception_pc_set                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.illegal_insn_q                                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.illegal_insn_q                                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.load_err_q                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.load_err_q                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.nmi_mode_q                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.nmi_mode_q                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.seen_exception_pc_set                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.seen_exception_pc_set                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.store_err_q                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.store_err_q                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.g_branch_set_flop.branch_set_raw_q                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.g_branch_set_flop.branch_set_raw_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.g_sec_branch_taken.branch_taken_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.g_sec_branch_taken.branch_taken_q                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.id_fsm_q                                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.id_fsm_q                                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.imd_val_q                                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.imd_val_q                                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.dummy_instr_id_o                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.dummy_instr_id_o                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.g_secure_pc.prev_instr_seq_q                                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.g_secure_pc.prev_instr_seq_q                                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_cnt_q                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_cnt_q                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_instr_seed_q                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_instr_seed_q                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.cnt_q                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.cnt_q                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.perturbed_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.perturbed_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.lfsr_q                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.lfsr_q                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_addr_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_addr_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_busy_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_busy_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_cache_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_cache_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_data_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_data_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_err_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_err_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_cnt_q                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_cnt_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_done_q                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_done_q                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_hold_q                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_hold_q                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_hit_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_hit_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_in_ic1                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_in_ic1                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_older_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_older_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_out_cnt_q                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_out_cnt_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ram_done_q                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ram_done_q                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_rvd_cnt_q                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_rvd_cnt_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_stale_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_stale_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_way_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_way_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_index_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_index_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_ways_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_ways_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_write_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_write_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.lookup_index_ic1                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.lookup_index_ic1                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.inval_index_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.inval_index_q                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.inval_prog_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.inval_prog_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.lookup_addr_ic1                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.lookup_addr_ic1                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.lookup_valid_ic1                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.lookup_valid_ic1                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.output_addr_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.output_addr_q                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.prefetch_addr_q                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.prefetch_addr_q                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.reset_inval_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.reset_inval_q                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.round_robin_way_q                                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.round_robin_way_q                                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_data_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_data_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_err_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_err_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_valid_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_valid_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.illegal_c_insn_id_o                                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.illegal_c_insn_id_o                                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_fetch_err_o                                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_fetch_err_o                                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_fetch_err_plus2_o                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_fetch_err_plus2_o                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_is_compressed_id_o                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_is_compressed_id_o                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_new_id_q                                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_new_id_q                                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_alu_id_o                                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_alu_id_o                                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_c_id_o                                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_c_id_o                                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_id_o                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_id_o                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_valid_id_q                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_valid_id_q                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.pc_id_o                                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.pc_id_o                                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.addr_last_q                                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.addr_last_q                                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_sign_ext_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_sign_ext_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_type_q                                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_type_q                                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_we_q                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_we_q                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.handle_misaligned_q                                                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.handle_misaligned_q                                                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.ls_fsm_cs                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.ls_fsm_cs                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.lsu_err_q                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.lsu_err_q                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.pmp_err_q                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.pmp_err_q                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.rdata_offset_q                                                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.rdata_offset_q                                                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.rdata_q                                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.rdata_q                                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_waddr_wb_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_waddr_wb_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_wdata_wb_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_wdata_wb_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_we_wb_q                                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_we_wb_q                                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_compressed_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_compressed_q                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_count_q                                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_count_q                                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_instr_type_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_instr_type_q                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_pc_q                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_pc_q                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_valid_q                                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_valid_q                                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_esc_receiver.state_q                                                                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_esc_receiver.state_q                                                                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_esc_receiver.u_decode_esc.gen_no_async.diff_pq                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_esc_receiver.u_decode_esc.gen_no_async.diff_pq                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_esc_receiver.u_decode_esc.level_q                                                                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_esc_receiver.u_decode_esc.level_q                                                                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_esc_receiver.u_prim_generic_flop.q_o                                                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_esc_receiver.u_prim_generic_flop.q_o                                                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_pwrmgr_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_pwrmgr_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_pwrmgr_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_pwrmgr_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o
    );
endfunction

function automatic soc_state_equivalence_rv_core_ibex();
    soc_state_equivalence_rv_core_ibex = (
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_d_ibex.g_multiple_reqs.source_q                                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_d_ibex.g_multiple_reqs.source_q                                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_d_ibex.intg_err_q                                                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_d_ibex.intg_err_q                                                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_d_ibex.outstanding_reqs_q                                                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_d_ibex.outstanding_reqs_q                                                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_i_ibex.g_multiple_reqs.source_q                                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_i_ibex.g_multiple_reqs.source_q                                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_i_ibex.intg_err_q                                                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_i_ibex.intg_err_q                                                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.tl_adapter_host_i_ibex.outstanding_reqs_q                                                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.tl_adapter_host_i_ibex.outstanding_reqs_q                                                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.core_busy_q                                                                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.core_busy_q                                                                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.core_clock_gate_i.gen_generic.u_impl_generic.en_latch                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.core_clock_gate_i.gen_generic.u_impl_generic.en_latch                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.fetch_enable_q                                                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.fetch_enable_q                                                                                                               &&
        //top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.core_outputs_q                                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.core_outputs_q                                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.rst_shadow_cnt_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.rst_shadow_cnt_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.rst_shadow_set_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.rst_shadow_set_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_data_rdata_q                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_data_rdata_q                                                                             &&
        //top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_inputs_q                                                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_inputs_q                                                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_tag_rdata_q                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.shadow_tag_rdata_q                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_addr_csr.rdata_q             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_addr_csr.rdata_q              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_cfg_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_cfg_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_addr_csr.rdata_q              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_addr_csr.rdata_q               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_cfg_csr.rdata_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_cfg_csr.rdata_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.u_pmp_mseccfg.rdata_q                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.g_pmp_registers.u_pmp_mseccfg.rdata_q                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[0].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[0].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[1].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[1].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[2].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[2].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[3].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[3].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[4].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[4].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[5].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[5].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[6].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[6].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[7].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[7].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[8].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[8].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[9].gen_imp.mcounters_variable_i.counter_q               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_cntrs[9].gen_imp.mcounters_variable_i.counter_q                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr.rdata_q == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr.rdata_q   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr.rdata_q    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.u_tselect_csr.rdata_q                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.gen_trigger_regs.u_tselect_csr.rdata_q                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.mcountinhibit_q                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.mcountinhibit_q                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.mcycle_counter_i.counter_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.mcycle_counter_i.counter_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.minstret_counter_i.counter_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.minstret_counter_i.counter_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.priv_lvl_q                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.priv_lvl_q                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_cpuctrl_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_cpuctrl_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dcsr_csr.rdata_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dcsr_csr.rdata_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_depc_csr.rdata_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_depc_csr.rdata_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dscratch0_csr.rdata_q                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dscratch0_csr.rdata_q                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dscratch1_csr.rdata_q                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_dscratch1_csr.rdata_q                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mcause_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mcause_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mepc_csr.rdata_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mepc_csr.rdata_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mie_csr.rdata_q                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mie_csr.rdata_q                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mscratch_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mscratch_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_cause_csr.rdata_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_cause_csr.rdata_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_epc_csr.rdata_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstack_epc_csr.rdata_q                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstatus_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mstatus_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mtval_csr.rdata_q                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mtval_csr.rdata_q                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mtvec_csr.rdata_q                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.cs_registers_i.u_mtvec_csr.rdata_q                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_single_cycle.mult_state_q         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_single_cycle.mult_state_q          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.branch_jump_set_done_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.branch_jump_set_done_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.ctrl_fsm_cs                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.ctrl_fsm_cs                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.debug_mode_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.debug_mode_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.do_single_step_q                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.do_single_step_q                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.enter_debug_mode_prio_q                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.enter_debug_mode_prio_q                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exc_req_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exc_req_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exception_req_accepted                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exception_req_accepted                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exception_req_pending                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.exception_req_pending                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.expect_exception_pc_set                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.expect_exception_pc_set                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.illegal_insn_q                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.illegal_insn_q                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.load_err_q                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.load_err_q                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.nmi_mode_q                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.nmi_mode_q                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.seen_exception_pc_set                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.seen_exception_pc_set                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.store_err_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.controller_i.store_err_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.g_branch_set_flop.branch_set_raw_q                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.g_branch_set_flop.branch_set_raw_q                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.g_sec_branch_taken.branch_taken_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.g_sec_branch_taken.branch_taken_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.id_fsm_q                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.id_fsm_q                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.imd_val_q                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.id_stage_i.imd_val_q                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.dummy_instr_id_o                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.dummy_instr_id_o                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.g_secure_pc.prev_instr_seq_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.g_secure_pc.prev_instr_seq_q                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_cnt_q                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_cnt_q                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_instr_seed_q                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_instr_seed_q                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.cnt_q            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.cnt_q             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.perturbed_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.perturbed_q       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.lfsr_q                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.lfsr_q                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_addr_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_addr_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_busy_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_busy_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_cache_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_cache_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_data_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_data_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_err_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_err_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_cnt_q                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_cnt_q                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_done_q                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_done_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_hold_q                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ext_hold_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_hit_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_hit_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_in_ic1                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_in_ic1                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_older_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_older_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_out_cnt_q                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_out_cnt_q                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ram_done_q                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_ram_done_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_rvd_cnt_q                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_rvd_cnt_q                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_stale_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_stale_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_way_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.fill_way_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_index_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_index_q       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_ways_q       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_ways_q        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_write_q      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_write_q       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.lookup_index_ic1            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.lookup_index_ic1             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.inval_index_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.inval_index_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.inval_prog_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.inval_prog_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.lookup_addr_ic1                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.lookup_addr_ic1                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.lookup_valid_ic1                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.lookup_valid_ic1                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.output_addr_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.output_addr_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.prefetch_addr_q                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.prefetch_addr_q                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.reset_inval_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.reset_inval_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.round_robin_way_q                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.round_robin_way_q                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_data_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_data_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_err_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_err_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_valid_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.gen_icache.icache_i.skid_valid_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.illegal_c_insn_id_o                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.illegal_c_insn_id_o                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_fetch_err_o                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_fetch_err_o                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_fetch_err_plus2_o                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_fetch_err_plus2_o                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_is_compressed_id_o                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_is_compressed_id_o                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_new_id_q                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_new_id_q                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_alu_id_o                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_alu_id_o                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_c_id_o                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_c_id_o                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_id_o                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_rdata_id_o                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_valid_id_q                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.instr_valid_id_q                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.pc_id_o                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.if_stage_i.pc_id_o                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.addr_last_q                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.addr_last_q                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_sign_ext_q                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_sign_ext_q                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_type_q                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_type_q                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_we_q                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.data_we_q                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.handle_misaligned_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.handle_misaligned_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.ls_fsm_cs                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.ls_fsm_cs                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.lsu_err_q                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.lsu_err_q                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.pmp_err_q                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.pmp_err_q                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.rdata_offset_q                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.rdata_offset_q                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.rdata_q                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.load_store_unit_i.rdata_q                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_waddr_wb_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_waddr_wb_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_wdata_wb_q                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_wdata_wb_q                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_we_wb_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.rf_we_wb_q                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_compressed_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_compressed_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_count_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_count_q                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_instr_type_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_instr_type_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_pc_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_pc_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_valid_q                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_lockstep.u_ibex_lockstep.u_shadow_core.wb_stage_i.g_writeback_stage.wb_valid_q                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].data_bank.gen_generic.u_impl_generic.mem                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].data_bank.gen_generic.u_impl_generic.mem                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].data_bank.gen_generic.u_impl_generic.rdata_o                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].data_bank.gen_generic.u_impl_generic.rdata_o                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].tag_bank.gen_generic.u_impl_generic.mem                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].tag_bank.gen_generic.u_impl_generic.mem                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].tag_bank.gen_generic.u_impl_generic.rdata_o                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[0].tag_bank.gen_generic.u_impl_generic.rdata_o                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].data_bank.gen_generic.u_impl_generic.mem                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].data_bank.gen_generic.u_impl_generic.mem                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].data_bank.gen_generic.u_impl_generic.rdata_o                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].data_bank.gen_generic.u_impl_generic.rdata_o                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].tag_bank.gen_generic.u_impl_generic.mem                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].tag_bank.gen_generic.u_impl_generic.mem                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].tag_bank.gen_generic.u_impl_generic.rdata_o                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_rams.gen_rams_inner[1].tag_bank.gen_generic.u_impl_generic.rdata_o                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_regfile_ff.register_file_i.g_dummy_r0.rf_r0_q                                                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_regfile_ff.register_file_i.g_dummy_r0.rf_r0_q                                                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.gen_regfile_ff.register_file_i.rf_reg_q                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.gen_regfile_ff.register_file_i.rf_reg_q                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[0].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[10].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[11].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[12].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[13].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[14].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_addr_csr.rdata_q                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_addr_csr.rdata_q                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_cfg_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[15].u_pmp_cfg_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[1].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[2].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[3].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[4].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[5].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[6].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[7].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[8].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_addr_csr.rdata_q                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_addr_csr.rdata_q                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_cfg_csr.rdata_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.g_pmp_csrs[9].u_pmp_cfg_csr.rdata_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.u_pmp_mseccfg.rdata_q                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.g_pmp_registers.u_pmp_mseccfg.rdata_q                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[0].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[0].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[1].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[1].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[2].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[2].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[3].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[3].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[4].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[4].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[5].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[5].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[6].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[6].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[7].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[7].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[8].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[8].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[9].gen_imp.mcounters_variable_i.counter_q                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_cntrs[9].gen_imp.mcounters_variable_i.counter_q                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr.rdata_q                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_control_csr.rdata_q                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr.rdata_q                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.g_dbg_tmatch_reg[0].u_tmatch_value_csr.rdata_q                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.u_tselect_csr.rdata_q                                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.gen_trigger_regs.u_tselect_csr.rdata_q                                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcountinhibit_q                                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcountinhibit_q                                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcycle_counter_i.counter_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.mcycle_counter_i.counter_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.minstret_counter_i.counter_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.minstret_counter_i.counter_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.priv_lvl_q                                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.priv_lvl_q                                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_cpuctrl_csr.rdata_q                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_cpuctrl_csr.rdata_q                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dcsr_csr.rdata_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dcsr_csr.rdata_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_depc_csr.rdata_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_depc_csr.rdata_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch0_csr.rdata_q                                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch0_csr.rdata_q                                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch1_csr.rdata_q                                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_dscratch1_csr.rdata_q                                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mcause_csr.rdata_q                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mcause_csr.rdata_q                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mepc_csr.rdata_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mepc_csr.rdata_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mie_csr.rdata_q                                                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mie_csr.rdata_q                                                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mscratch_csr.rdata_q                                                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mscratch_csr.rdata_q                                                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_cause_csr.rdata_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_cause_csr.rdata_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_csr.rdata_q                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_csr.rdata_q                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_epc_csr.rdata_q                                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstack_epc_csr.rdata_q                                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstatus_csr.rdata_q                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mstatus_csr.rdata_q                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtval_csr.rdata_q                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtval_csr.rdata_q                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtvec_csr.rdata_q                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.cs_registers_i.u_mtvec_csr.rdata_q                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_single_cycle.mult_state_q                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_single_cycle.mult_state_q                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q                                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q                                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.branch_jump_set_done_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.branch_jump_set_done_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.ctrl_fsm_cs                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.ctrl_fsm_cs                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.debug_mode_q                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.debug_mode_q                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.do_single_step_q                                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.do_single_step_q                                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.enter_debug_mode_prio_q                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.enter_debug_mode_prio_q                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exc_req_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exc_req_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exception_req_accepted                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exception_req_accepted                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exception_req_pending                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.exception_req_pending                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.expect_exception_pc_set                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.expect_exception_pc_set                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.illegal_insn_q                                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.illegal_insn_q                                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.load_err_q                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.load_err_q                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.nmi_mode_q                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.nmi_mode_q                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.seen_exception_pc_set                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.seen_exception_pc_set                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.store_err_q                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.controller_i.store_err_q                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.g_branch_set_flop.branch_set_raw_q                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.g_branch_set_flop.branch_set_raw_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.g_sec_branch_taken.branch_taken_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.g_sec_branch_taken.branch_taken_q                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.id_fsm_q                                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.id_fsm_q                                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.imd_val_q                                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.id_stage_i.imd_val_q                                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.dummy_instr_id_o                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.dummy_instr_id_o                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.g_secure_pc.prev_instr_seq_q                                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.g_secure_pc.prev_instr_seq_q                                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_cnt_q                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_cnt_q                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_instr_seed_q                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_instr_seed_q                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.cnt_q                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.cnt_q                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.perturbed_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.gen_max_len_sva.perturbed_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.lfsr_q                                                          == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_i.lfsr_q                                                           &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_addr_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_addr_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_busy_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_busy_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_cache_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_cache_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_data_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_data_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_err_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_err_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_cnt_q                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_cnt_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_done_q                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_done_q                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_hold_q                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ext_hold_q                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_hit_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_hit_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_in_ic1                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_in_ic1                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_older_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_older_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_out_cnt_q                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_out_cnt_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ram_done_q                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_ram_done_q                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_rvd_cnt_q                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_rvd_cnt_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_stale_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_stale_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_way_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.fill_way_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_index_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_index_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_ways_q                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_ways_q                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_write_q                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.ecc_correction_write_q                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.lookup_index_ic1                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.gen_data_ecc_checking.lookup_index_ic1                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.inval_index_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.inval_index_q                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.inval_prog_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.inval_prog_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.lookup_addr_ic1                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.lookup_addr_ic1                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.lookup_valid_ic1                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.lookup_valid_ic1                                                                  &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.output_addr_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.output_addr_q                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.prefetch_addr_q                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.prefetch_addr_q                                                                   &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.reset_inval_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.reset_inval_q                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.round_robin_way_q                                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.round_robin_way_q                                                                 &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_data_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_data_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_err_q                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_err_q                                                                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_valid_q                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.gen_icache.icache_i.skid_valid_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.illegal_c_insn_id_o                                                                                  == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.illegal_c_insn_id_o                                                                                   &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_fetch_err_o                                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_fetch_err_o                                                                                     &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_fetch_err_plus2_o                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_fetch_err_plus2_o                                                                               &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_is_compressed_id_o                                                                             == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_is_compressed_id_o                                                                              &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_new_id_q                                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_new_id_q                                                                                        &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_alu_id_o                                                                                 == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_alu_id_o                                                                                  &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_c_id_o                                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_c_id_o                                                                                    &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_id_o                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_rdata_id_o                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_valid_id_q                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.instr_valid_id_q                                                                                      &&
 //       top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.pc_id_o                                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.if_stage_i.pc_id_o                                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.addr_last_q                                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.addr_last_q                                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_sign_ext_q                                                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_sign_ext_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_type_q                                                                                   == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_type_q                                                                                    &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_we_q                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.data_we_q                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.handle_misaligned_q                                                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.handle_misaligned_q                                                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.ls_fsm_cs                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.ls_fsm_cs                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.lsu_err_q                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.lsu_err_q                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.pmp_err_q                                                                                     == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.pmp_err_q                                                                                      &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.rdata_offset_q                                                                                == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.rdata_offset_q                                                                                 &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.rdata_q                                                                                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.load_store_unit_i.rdata_q                                                                                        &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_waddr_wb_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_waddr_wb_q                                                                       &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_wdata_wb_q                                                                      == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_wdata_wb_q                                                                       &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_we_wb_q                                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.rf_we_wb_q                                                                          &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_compressed_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_compressed_q                                                                     &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_count_q                                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_count_q                                                                          &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_instr_type_q                                                                    == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_instr_type_q                                                                     &&
//        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_pc_q                                                                            == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_pc_q                                                                             &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_valid_q                                                                         == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_core.u_ibex_core.wb_stage_i.g_writeback_stage.wb_valid_q                                                                          &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_esc_receiver.state_q                                                                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_esc_receiver.state_q                                                                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_esc_receiver.u_decode_esc.gen_no_async.diff_pq                                                                              == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_esc_receiver.u_decode_esc.gen_no_async.diff_pq                                                                               &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_esc_receiver.u_decode_esc.level_q                                                                                           == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_esc_receiver.u_decode_esc.level_q                                                                                            &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_esc_receiver.u_prim_generic_flop.q_o                                                                                        == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_esc_receiver.u_prim_generic_flop.q_o                                                                                         &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                                               == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                                                &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_pwrmgr_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_pwrmgr_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                        &&
        top_level_upec.top_earlgrey_1.u_rv_core_ibex.u_pwrmgr_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_rv_core_ibex.u_pwrmgr_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o
    );
endfunction