function automatic black_box_input_equivalence_peri_devices();
    black_box_input_equivalence_peri_devices = (
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.rdata_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.rdata_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o                                       == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o                                    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o                                       == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o                                    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o                                           == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o                                        &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o                                           == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o
        );
endfunction

function automatic black_box_output_equivalence_peri_devices();
    black_box_output_equivalence_peri_devices = (
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.addr_i     == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.addr_i  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.cfg_i      == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.addr_i  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.clk_i      == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.addr_i  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.req_i      == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.addr_i  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.wdata_i    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.addr_i  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.wmask_i    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.addr_i  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.write_i    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.addr_i  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_addr_i                                        == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_addr_i                                     &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_req_i                                         == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_req_i                                      &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_wdata_i                                       == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_wdata_i                                    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_wmask_i                                       == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_wmask_i                                    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_write_i                                       == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_write_i                                    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_addr_i                                        == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_addr_i                                     &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_req_i                                         == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_req_i                                      &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_wdata_i                                       == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_wdata_i                                    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_wmask_i                                       == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_wmask_i                                    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_write_i                                       == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_write_i                                    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.cfg_i                                           == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.cfg_i                                        &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.clk_a_i                                         == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.clk_a_i                                      &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.clk_b_i                                         == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.clk_b_i                                      &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_addr_i                                            == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_addr_i                                         &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_req_i                                             == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_req_i                                          &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_wdata_i                                           == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_wdata_i                                        &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_wmask_i                                           == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_wmask_i                                        &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_write_i                                           == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_write_i                                        &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_addr_i                                            == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_addr_i                                         &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_req_i                                             == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_req_i                                          &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_wdata_i                                           == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_wdata_i                                        &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_wmask_i                                           == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_wmask_i                                        &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_write_i                                           == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_write_i                                        &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.cfg_i                                               == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.cfg_i                                            &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.clk_a_i                                             == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.clk_a_i                                          &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.clk_b_i                                             == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.clk_b_i
    );
endfunction

function automatic input_equivalence_peri_devices();
    input_equivalence_peri_devices = (
//        top_level_upec.top_earlgrey_1.u_uart0.cio_rx_i      == top_level_upec.top_earlgrey_2.u_uart0.cio_rx_i   && 
//        top_level_upec.top_earlgrey_1.u_uart0.alert_rx_i    == top_level_upec.top_earlgrey_2.u_uart0.alert_rx_i && 
//        top_level_upec.top_earlgrey_1.u_uart0.tl_i          == top_level_upec.top_earlgrey_2.u_uart0.tl_i       && 
//        top_level_upec.top_earlgrey_1.u_uart0.clk_i         == top_level_upec.top_earlgrey_2.u_uart0.clk_i      && 
//        top_level_upec.top_earlgrey_1.u_uart0.rst_ni        == top_level_upec.top_earlgrey_2.u_uart0.rst_ni     &&

//        top_level_upec.top_earlgrey_1.u_uart1.cio_rx_i      == top_level_upec.top_earlgrey_2.u_uart1.cio_rx_i   && 
//        top_level_upec.top_earlgrey_1.u_uart1.alert_rx_i    == top_level_upec.top_earlgrey_2.u_uart1.alert_rx_i && 
//        top_level_upec.top_earlgrey_1.u_uart1.tl_i          == top_level_upec.top_earlgrey_2.u_uart1.tl_i       && 
//        top_level_upec.top_earlgrey_1.u_uart1.clk_i         == top_level_upec.top_earlgrey_2.u_uart1.clk_i      && 
//        top_level_upec.top_earlgrey_1.u_uart1.rst_ni        == top_level_upec.top_earlgrey_2.u_uart1.rst_ni     &&

//        top_level_upec.top_earlgrey_1.u_uart2.cio_rx_i      == top_level_upec.top_earlgrey_2.u_uart2.cio_rx_i   && 
//        top_level_upec.top_earlgrey_1.u_uart2.alert_rx_i    == top_level_upec.top_earlgrey_2.u_uart2.alert_rx_i && 
//        top_level_upec.top_earlgrey_1.u_uart2.tl_i          == top_level_upec.top_earlgrey_2.u_uart2.tl_i       && 
//        top_level_upec.top_earlgrey_1.u_uart2.clk_i         == top_level_upec.top_earlgrey_2.u_uart2.clk_i      && 
//        top_level_upec.top_earlgrey_1.u_uart2.rst_ni        == top_level_upec.top_earlgrey_2.u_uart2.rst_ni     &&

//        top_level_upec.top_earlgrey_1.u_uart3.cio_rx_i      == top_level_upec.top_earlgrey_2.u_uart3.cio_rx_i   && 
//        top_level_upec.top_earlgrey_1.u_uart3.alert_rx_i    == top_level_upec.top_earlgrey_2.u_uart3.alert_rx_i && 
//        top_level_upec.top_earlgrey_1.u_uart3.tl_i          == top_level_upec.top_earlgrey_2.u_uart3.tl_i       && 
//        top_level_upec.top_earlgrey_1.u_uart3.clk_i         == top_level_upec.top_earlgrey_2.u_uart3.clk_i      && 
//        top_level_upec.top_earlgrey_1.u_uart3.rst_ni        == top_level_upec.top_earlgrey_2.u_uart3.rst_ni     && 

//        top_level_upec.top_earlgrey_1.u_spi_host0.cio_sd_i  == top_level_upec.top_earlgrey_2.u_spi_host0.cio_sd_i   &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.alert_rx_i    == top_level_upec.top_earlgrey_2.u_spi_host0.alert_rx_i &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.passthrough_i == top_level_upec.top_earlgrey_2.u_spi_host0.passthrough_i  &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.tl_i  == top_level_upec.top_earlgrey_2.u_spi_host0.tl_i   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.scanmode_i    == top_level_upec.top_earlgrey_2.u_spi_host0.scanmode_i &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.clk_i == top_level_upec.top_earlgrey_2.u_spi_host0.clk_i  &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.clk_core_i    == top_level_upec.top_earlgrey_2.u_spi_host0.clk_core_i &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.rst_ni    == top_level_upec.top_earlgrey_2.u_spi_host0.rst_ni &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.rst_core_ni   == top_level_upec.top_earlgrey_2.u_spi_host0.rst_core_ni    &&

//        top_level_upec.top_earlgrey_1.u_spi_host1.cio_sd_i  == top_level_upec.top_earlgrey_2.u_spi_host1.cio_sd_i   &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.alert_rx_i    == top_level_upec.top_earlgrey_2.u_spi_host1.alert_rx_i &&
        top_level_upec.top_earlgrey_1.u_spi_host1.passthrough_i == top_level_upec.top_earlgrey_2.u_spi_host1.passthrough_i  &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.tl_i  == top_level_upec.top_earlgrey_2.u_spi_host1.tl_i   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.scanmode_i    == top_level_upec.top_earlgrey_2.u_spi_host1.scanmode_i &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.clk_i == top_level_upec.top_earlgrey_2.u_spi_host1.clk_i  &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.clk_core_i    == top_level_upec.top_earlgrey_2.u_spi_host1.clk_core_i &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.rst_ni    == top_level_upec.top_earlgrey_2.u_spi_host1.rst_ni &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.rst_core_ni   == top_level_upec.top_earlgrey_2.u_spi_host1.rst_core_ni    &&

//        top_level_upec.top_earlgrey_1.u_spi_device.cio_sck_i    == top_level_upec.top_earlgrey_2.u_spi_device.cio_sck_i &&
//        top_level_upec.top_earlgrey_1.u_spi_device.cio_csb_i    == top_level_upec.top_earlgrey_2.u_spi_device.cio_csb_i &&
//        top_level_upec.top_earlgrey_1.u_spi_device.cio_sd_i == top_level_upec.top_earlgrey_2.u_spi_device.cio_sd_i  &&
//        top_level_upec.top_earlgrey_1.u_spi_device.alert_rx_i   == top_level_upec.top_earlgrey_2.u_spi_device.alert_rx_i    &&
        top_level_upec.top_earlgrey_1.u_spi_device.ram_cfg_i    == top_level_upec.top_earlgrey_2.u_spi_device.ram_cfg_i &&
//        top_level_upec.top_earlgrey_1.u_spi_device.passthrough_i    == top_level_upec.top_earlgrey_2.u_spi_device.passthrough_i &&
        top_level_upec.top_earlgrey_1.u_spi_device.mbist_en_i   == top_level_upec.top_earlgrey_2.u_spi_device.mbist_en_i    &&
//        top_level_upec.top_earlgrey_1.u_spi_device.tl_i == top_level_upec.top_earlgrey_2.u_spi_device.tl_i  &&
        top_level_upec.top_earlgrey_1.u_spi_device.scanmode_i   == top_level_upec.top_earlgrey_2.u_spi_device.scanmode_i    &&
        top_level_upec.top_earlgrey_1.u_spi_device.scan_rst_ni  == top_level_upec.top_earlgrey_2.u_spi_device.scan_rst_ni   &&
//        top_level_upec.top_earlgrey_1.u_spi_device.clk_i    == top_level_upec.top_earlgrey_2.u_spi_device.clk_i &&
//        top_level_upec.top_earlgrey_1.u_spi_device.scan_clk_i   == top_level_upec.top_earlgrey_2.u_spi_device.scan_clk_i    &&
//        top_level_upec.top_earlgrey_1.u_spi_device.rst_ni   == top_level_upec.top_earlgrey_2.u_spi_device.rst_ni    &&

//        top_level_upec.top_earlgrey_1.u_usbdev.cio_sense_i   == top_level_upec.top_earlgrey_2.u_usbdev.cio_sense_i    &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_d_i   == top_level_upec.top_earlgrey_2.u_usbdev.cio_d_i    &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_dp_i  == top_level_upec.top_earlgrey_2.u_usbdev.cio_dp_i   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_dn_i  == top_level_upec.top_earlgrey_2.u_usbdev.cio_dn_i   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.usb_state_debug_i == top_level_upec.top_earlgrey_2.u_usbdev.usb_state_debug_i  &&
        top_level_upec.top_earlgrey_1.u_usbdev.ram_cfg_i == top_level_upec.top_earlgrey_2.u_usbdev.ram_cfg_i  &&
//        top_level_upec.top_earlgrey_1.u_usbdev.tl_i  == top_level_upec.top_earlgrey_2.u_usbdev.tl_i   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.clk_i == top_level_upec.top_earlgrey_2.u_usbdev.clk_i  &&
//        top_level_upec.top_earlgrey_1.u_usbdev.clk_aon_i == top_level_upec.top_earlgrey_2.u_usbdev.clk_aon_i  &&
//        top_level_upec.top_earlgrey_1.u_usbdev.clk_usb_48mhz_i   == top_level_upec.top_earlgrey_2.u_usbdev.clk_usb_48mhz_i    &&
//        top_level_upec.top_earlgrey_1.u_usbdev.rst_ni    == top_level_upec.top_earlgrey_2.u_usbdev.rst_ni &&
//        top_level_upec.top_earlgrey_1.u_usbdev.rst_aon_ni    == top_level_upec.top_earlgrey_2.u_usbdev.rst_aon_ni &&
//        top_level_upec.top_earlgrey_1.u_usbdev.rst_usb_48mhz_ni  == top_level_upec.top_earlgrey_2.u_usbdev.rst_usb_48mhz_ni   &&

//        top_level_upec.top_earlgrey_1.u_gpio.cio_gpio_i == top_level_upec.top_earlgrey_2.u_gpio.cio_gpio_i  &&
//        top_level_upec.top_earlgrey_1.u_gpio.alert_rx_i == top_level_upec.top_earlgrey_2.u_gpio.alert_rx_i  &&
//        top_level_upec.top_earlgrey_1.u_gpio.tl_i   == top_level_upec.top_earlgrey_2.u_gpio.tl_i    &&
//        top_level_upec.top_earlgrey_1.u_gpio.clk_i  == top_level_upec.top_earlgrey_2.u_gpio.clk_i   &&
//        top_level_upec.top_earlgrey_1.u_gpio.rst_ni == top_level_upec.top_earlgrey_2.u_gpio.rst_ni  &&

//        top_level_upec.top_earlgrey_1.u_i2c0.cio_sda_i  == top_level_upec.top_earlgrey_2.u_i2c0.cio_sda_i   &&
//        top_level_upec.top_earlgrey_1.u_i2c0.cio_scl_i  == top_level_upec.top_earlgrey_2.u_i2c0.cio_scl_i   &&
//        top_level_upec.top_earlgrey_1.u_i2c0.alert_rx_i == top_level_upec.top_earlgrey_2.u_i2c0.alert_rx_i  &&
//        top_level_upec.top_earlgrey_1.u_i2c0.tl_i   == top_level_upec.top_earlgrey_2.u_i2c0.tl_i    &&
//        top_level_upec.top_earlgrey_1.u_i2c0.clk_i  == top_level_upec.top_earlgrey_2.u_i2c0.clk_i   &&
//        top_level_upec.top_earlgrey_1.u_i2c0.rst_ni == top_level_upec.top_earlgrey_2.u_i2c0.rst_ni  &&

//        top_level_upec.top_earlgrey_1.u_i2c1.cio_sda_i  == top_level_upec.top_earlgrey_2.u_i2c1.cio_sda_i   &&
//        top_level_upec.top_earlgrey_1.u_i2c1.cio_scl_i  == top_level_upec.top_earlgrey_2.u_i2c1.cio_scl_i   &&
//        top_level_upec.top_earlgrey_1.u_i2c1.alert_rx_i == top_level_upec.top_earlgrey_2.u_i2c1.alert_rx_i  &&
//        top_level_upec.top_earlgrey_1.u_i2c1.tl_i   == top_level_upec.top_earlgrey_2.u_i2c1.tl_i    &&
//        top_level_upec.top_earlgrey_1.u_i2c1.clk_i  == top_level_upec.top_earlgrey_2.u_i2c1.clk_i   &&
//        top_level_upec.top_earlgrey_1.u_i2c1.rst_ni == top_level_upec.top_earlgrey_2.u_i2c1.rst_ni  &&

//        top_level_upec.top_earlgrey_1.u_i2c2.cio_sda_i  == top_level_upec.top_earlgrey_2.u_i2c2.cio_sda_i   &&
//        top_level_upec.top_earlgrey_1.u_i2c2.cio_scl_i  == top_level_upec.top_earlgrey_2.u_i2c2.cio_scl_i   &&
//        top_level_upec.top_earlgrey_1.u_i2c2.alert_rx_i == top_level_upec.top_earlgrey_2.u_i2c2.alert_rx_i  &&
//        top_level_upec.top_earlgrey_1.u_i2c2.tl_i   == top_level_upec.top_earlgrey_2.u_i2c2.tl_i    &&
//        top_level_upec.top_earlgrey_1.u_i2c2.clk_i  == top_level_upec.top_earlgrey_2.u_i2c2.clk_i   &&
//        top_level_upec.top_earlgrey_1.u_i2c2.rst_ni == top_level_upec.top_earlgrey_2.u_i2c2.rst_ni  &&

//        top_level_upec.top_earlgrey_1.u_pwm_aon.tl_i    == top_level_upec.top_earlgrey_2.u_pwm_aon.tl_i &&
//        top_level_upec.top_earlgrey_1.u_pwm_aon.clk_i   == top_level_upec.top_earlgrey_2.u_pwm_aon.clk_i    &&
//        top_level_upec.top_earlgrey_1.u_pwm_aon.clk_core_i  == top_level_upec.top_earlgrey_2.u_pwm_aon.clk_core_i   &&
//        top_level_upec.top_earlgrey_1.u_pwm_aon.rst_ni  == top_level_upec.top_earlgrey_2.u_pwm_aon.rst_ni   &&
//        top_level_upec.top_earlgrey_1.u_pwm_aon.rst_core_ni == top_level_upec.top_earlgrey_2.u_pwm_aon.rst_core_ni  &&


//        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.alert_rx_i == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.alert_rx_i  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.adc_i  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.adc_i   &&
//        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.tl_i   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.tl_i    &&
//        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.clk_i  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.clk_i   &&
//        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.clk_aon_i  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.clk_aon_i   &&
//        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.rst_ni == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.rst_ni  &&
//        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.rst_slow_ni    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.rst_slow_ni &&

//        top_level_upec.top_earlgrey_1.u_rstmgr_aon.pwr_i    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.pwr_i &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.cpu_i    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.cpu_i &&
//        top_level_upec.top_earlgrey_1.u_rstmgr_aon.alert_dump_i == top_level_upec.top_earlgrey_2.u_rstmgr_aon.alert_dump_i  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.cpu_dump_i   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.cpu_dump_i    &&
//        top_level_upec.top_earlgrey_1.u_rstmgr_aon.tl_i == top_level_upec.top_earlgrey_2.u_rstmgr_aon.tl_i  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.scanmode_i   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.scanmode_i    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.scan_rst_ni  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.scan_rst_ni   &&
//        top_level_upec.top_earlgrey_1.u_rstmgr_aon.clk_i    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.clk_i &&
//        top_level_upec.top_earlgrey_1.u_rstmgr_aon.clk_aon_i    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.clk_aon_i &&
//        top_level_upec.top_earlgrey_1.u_rstmgr_aon.clk_main_i   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.clk_main_i    &&
//        top_level_upec.top_earlgrey_1.u_rstmgr_aon.clk_io_i == top_level_upec.top_earlgrey_2.u_rstmgr_aon.clk_io_i  &&
//        top_level_upec.top_earlgrey_1.u_rstmgr_aon.clk_usb_i    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.clk_usb_i &&
//        top_level_upec.top_earlgrey_1.u_rstmgr_aon.clk_io_div2_i    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.clk_io_div2_i &&
//        top_level_upec.top_earlgrey_1.u_rstmgr_aon.clk_io_div4_i    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.clk_io_div4_i &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.rst_ni   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.rst_ni    &&

//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.lc_dft_en_i  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.lc_dft_en_i   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.ast_clk_byp_ack_i    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.ast_clk_byp_ack_i &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.lc_clk_byp_req_i == top_level_upec.top_earlgrey_2.u_clkmgr_aon.lc_clk_byp_req_i  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.clk_main_i   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.clk_main_i    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.clk_io_i == top_level_upec.top_earlgrey_2.u_clkmgr_aon.clk_io_i  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.clk_usb_i    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.clk_usb_i &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.clk_aon_i    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.clk_aon_i &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.pwr_i    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.pwr_i &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.idle_i   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.idle_i    &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.tl_i == top_level_upec.top_earlgrey_2.u_clkmgr_aon.tl_i  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.scanmode_i   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.scanmode_i    &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.clk_i    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.clk_i &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.rst_ni   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.rst_ni    &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.rst_main_ni  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.rst_main_ni   &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.rst_io_ni    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.rst_io_ni &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.rst_usb_ni   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.rst_usb_ni    &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.rst_io_div2_ni   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.rst_io_div2_ni    &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.rst_io_div4_ni   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.rst_io_div4_ni    &&

        
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_ast_i    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_ast_i &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_rst_i    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_rst_i &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_clk_i    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_clk_i &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_otp_i    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_otp_i &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_lc_i == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_lc_i  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_flash_i  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_flash_i   &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.esc_rst_tx_i == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.esc_rst_tx_i  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_cpu_i    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_cpu_i &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.wakeups_i    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.wakeups_i &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.rstreqs_i    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.rstreqs_i &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.rom_ctrl_i   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.rom_ctrl_i    &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.tl_i == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.tl_i  &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.clk_i    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.clk_i &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.clk_slow_i   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.clk_slow_i    &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.rst_ni   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.rst_ni    &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.rst_slow_ni  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.rst_slow_ni   &&

//        top_level_upec.top_earlgrey_1.u_rv_timer.tl_i   == top_level_upec.top_earlgrey_2.u_rv_timer.tl_i    &&
//        top_level_upec.top_earlgrey_1.u_rv_timer.clk_i  == top_level_upec.top_earlgrey_2.u_rv_timer.clk_i   &&
//        top_level_upec.top_earlgrey_1.u_rv_timer.rst_ni == top_level_upec.top_earlgrey_2.u_rv_timer.rst_ni  &&

        top_level_upec.top_earlgrey_1.u_alert_handler.edn_i == top_level_upec.top_earlgrey_2.u_alert_handler.edn_i  &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.esc_rx_i  == top_level_upec.top_earlgrey_2.u_alert_handler.esc_rx_i   &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.tl_i  == top_level_upec.top_earlgrey_2.u_alert_handler.tl_i   &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.alert_tx_i[31:0]    == top_level_upec.top_earlgrey_2.u_alert_handler.alert_tx_i[31:0] &&
        top_level_upec.top_earlgrey_1.u_alert_handler.alert_tx_i[51:32]    == top_level_upec.top_earlgrey_2.u_alert_handler.alert_tx_i[51:32] &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.clk_i == top_level_upec.top_earlgrey_2.u_alert_handler.clk_i  &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.clk_edn_i == top_level_upec.top_earlgrey_2.u_alert_handler.clk_edn_i  &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.rst_ni    == top_level_upec.top_earlgrey_2.u_alert_handler.rst_ni &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.rst_edn_ni    == top_level_upec.top_earlgrey_2.u_alert_handler.rst_edn_ni &&

//        top_level_upec.top_earlgrey_1.u_aon_timer_aon.lc_escalate_en_i  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.lc_escalate_en_i   &&
//        top_level_upec.top_earlgrey_1.u_aon_timer_aon.sleep_mode_i  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.sleep_mode_i   &&
//        top_level_upec.top_earlgrey_1.u_aon_timer_aon.tl_i  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.tl_i   &&
//        top_level_upec.top_earlgrey_1.u_aon_timer_aon.clk_i == top_level_upec.top_earlgrey_2.u_aon_timer_aon.clk_i  &&
//        top_level_upec.top_earlgrey_1.u_aon_timer_aon.clk_aon_i == top_level_upec.top_earlgrey_2.u_aon_timer_aon.clk_aon_i  &&
//        top_level_upec.top_earlgrey_1.u_aon_timer_aon.rst_ni    == top_level_upec.top_earlgrey_2.u_aon_timer_aon.rst_ni &&
//        top_level_upec.top_earlgrey_1.u_aon_timer_aon.rst_aon_ni    == top_level_upec.top_earlgrey_2.u_aon_timer_aon.rst_aon_ni &&

//        top_level_upec.top_earlgrey_1.u_otp_ctrl.alert_rx_i == top_level_upec.top_earlgrey_2.u_otp_ctrl.alert_rx_i  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.otp_ast_pwr_seq_h_i    == top_level_upec.top_earlgrey_2.u_otp_ctrl.otp_ast_pwr_seq_h_i &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.edn_i  == top_level_upec.top_earlgrey_2.u_otp_ctrl.edn_i   &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.pwr_otp_i  == top_level_upec.top_earlgrey_2.u_otp_ctrl.pwr_otp_i   &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.lc_otp_program_i   == top_level_upec.top_earlgrey_2.u_otp_ctrl.lc_otp_program_i    &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.lc_escalate_en_i   == top_level_upec.top_earlgrey_2.u_otp_ctrl.lc_escalate_en_i    &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.lc_creator_seed_sw_rw_en_i == top_level_upec.top_earlgrey_2.u_otp_ctrl.lc_creator_seed_sw_rw_en_i  &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.lc_seed_hw_rd_en_i == top_level_upec.top_earlgrey_2.u_otp_ctrl.lc_seed_hw_rd_en_i  &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.lc_dft_en_i    == top_level_upec.top_earlgrey_2.u_otp_ctrl.lc_dft_en_i &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.lc_check_byp_en_i  == top_level_upec.top_earlgrey_2.u_otp_ctrl.lc_check_byp_en_i   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.flash_otp_key_i    == top_level_upec.top_earlgrey_2.u_otp_ctrl.flash_otp_key_i &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.sram_otp_key_i[0] == top_level_upec.top_earlgrey_2.u_otp_ctrl.sram_otp_key_i[0]  &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.sram_otp_key_i[1] == top_level_upec.top_earlgrey_2.u_otp_ctrl.sram_otp_key_i[1]  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.otbn_otp_key_i == top_level_upec.top_earlgrey_2.u_otp_ctrl.otbn_otp_key_i  &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.tl_i   == top_level_upec.top_earlgrey_2.u_otp_ctrl.tl_i    &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.otp_ext_voltage_h_io   == top_level_upec.top_earlgrey_2.u_otp_ctrl.otp_ext_voltage_h_io    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.scanmode_i == top_level_upec.top_earlgrey_2.u_otp_ctrl.scanmode_i  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.scan_rst_ni    == top_level_upec.top_earlgrey_2.u_otp_ctrl.scan_rst_ni &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.scan_en_i  == top_level_upec.top_earlgrey_2.u_otp_ctrl.scan_en_i   &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.clk_i  == top_level_upec.top_earlgrey_2.u_otp_ctrl.clk_i   &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.clk_edn_i  == top_level_upec.top_earlgrey_2.u_otp_ctrl.clk_edn_i   &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.rst_ni == top_level_upec.top_earlgrey_2.u_otp_ctrl.rst_ni  &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.rst_edn_ni == top_level_upec.top_earlgrey_2.u_otp_ctrl.rst_edn_ni  &&

//        top_level_upec.top_earlgrey_1.u_lc_ctrl.alert_rx_i    == top_level_upec.top_earlgrey_2.u_lc_ctrl.alert_rx_i &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.jtag_i    == top_level_upec.top_earlgrey_2.u_lc_ctrl.jtag_i &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.esc_wipe_secrets_tx_i == top_level_upec.top_earlgrey_2.u_lc_ctrl.esc_wipe_secrets_tx_i  &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.esc_scrap_state_tx_i  == top_level_upec.top_earlgrey_2.u_lc_ctrl.esc_scrap_state_tx_i   &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.pwr_lc_i  == top_level_upec.top_earlgrey_2.u_lc_ctrl.pwr_lc_i   &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.otp_lc_data_i == top_level_upec.top_earlgrey_2.u_lc_ctrl.otp_lc_data_i  &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_otp_program_i  == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_otp_program_i   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.kmac_data_i   == top_level_upec.top_earlgrey_2.u_lc_ctrl.kmac_data_i    &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_clk_byp_ack_i  == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_clk_byp_ack_i   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_flash_rma_ack_i    == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_flash_rma_ack_i &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.otp_device_id_i   == top_level_upec.top_earlgrey_2.u_lc_ctrl.otp_device_id_i    &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.tl_i  == top_level_upec.top_earlgrey_2.u_lc_ctrl.tl_i   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.scanmode_i    == top_level_upec.top_earlgrey_2.u_lc_ctrl.scanmode_i &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.scan_rst_ni   == top_level_upec.top_earlgrey_2.u_lc_ctrl.scan_rst_ni    &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.clk_i == top_level_upec.top_earlgrey_2.u_lc_ctrl.clk_i  &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.clk_kmac_i    == top_level_upec.top_earlgrey_2.u_lc_ctrl.clk_kmac_i &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.rst_ni    == top_level_upec.top_earlgrey_2.u_lc_ctrl.rst_ni &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.rst_kmac_ni   == top_level_upec.top_earlgrey_2.u_lc_ctrl.rst_kmac_ni    &&

//        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.clk_i    == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.clk_i &&
//        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.rst_ni   == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.rst_ni    &&
//        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.tl_i == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.tl_i  &&
//        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.en_ifetch_i  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.en_ifetch_i   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.gnt_i    == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.gnt_i &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.rdata_i  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.rdata_i   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.rvalid_i == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.rvalid_i  &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.rerror_i == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.rerror_i  &&

//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.alert_rx_i    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.alert_rx_i &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.sram_otp_key_i    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.sram_otp_key_i &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.sram_scr_i    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.sram_scr_i &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.sram_scr_init_i   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.sram_scr_init_i    &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.lc_escalate_en_i  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.lc_escalate_en_i   &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.lc_hw_debug_en_i  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.lc_hw_debug_en_i   &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.otp_en_sram_ifetch_i  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.otp_en_sram_ifetch_i   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.intg_error_i  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.intg_error_i   &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.tl_i  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.tl_i   &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.clk_i == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.clk_i  &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.clk_otp_i == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.clk_otp_i  &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.rst_ni    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.rst_ni &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.rst_otp_ni    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.rst_otp_ni &&

//        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.alert_rx_i  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.alert_rx_i   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.ast_alert_i == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.ast_alert_i  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.ast_status_i    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.ast_status_i &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.ast_init_done_i == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.ast_init_done_i  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.ast2pinmux_i    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.ast2pinmux_i &&
//        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.tl_i    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.tl_i &&
//        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.clk_i   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.clk_i    &&
//        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.rst_ni  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.rst_ni   &&

//        top_level_upec.top_earlgrey_1.u_pattgen.alert_rx_i  == top_level_upec.top_earlgrey_2.u_pattgen.alert_rx_i   &&
//        top_level_upec.top_earlgrey_1.u_pattgen.tl_i    == top_level_upec.top_earlgrey_2.u_pattgen.tl_i &&
//        top_level_upec.top_earlgrey_1.u_pattgen.clk_i   == top_level_upec.top_earlgrey_2.u_pattgen.clk_i    &&
//        top_level_upec.top_earlgrey_1.u_pattgen.rst_ni  == top_level_upec.top_earlgrey_2.u_pattgen.rst_ni   &&

//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_ac_present_i    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_ac_present_i &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_ec_rst_in_l_i   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_ec_rst_in_l_i    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_key0_in_i   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_key0_in_i    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_key1_in_i   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_key1_in_i    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_key2_in_i   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_key2_in_i    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_pwrb_in_i   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_pwrb_in_i    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.tl_i    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.tl_i &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.clk_i   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.clk_i    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.clk_aon_i   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.clk_aon_i    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.rst_ni  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.rst_ni   &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.rst_aon_ni  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.rst_aon_ni   &&

//        top_level_upec.top_earlgrey_1.u_pinmux_aon.alert_rx_i   == top_level_upec.top_earlgrey_2.u_pinmux_aon.alert_rx_i    &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.lc_hw_debug_en_i == top_level_upec.top_earlgrey_2.u_pinmux_aon.lc_hw_debug_en_i  &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.lc_dft_en_i  == top_level_upec.top_earlgrey_2.u_pinmux_aon.lc_dft_en_i   &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.lc_jtag_i    == top_level_upec.top_earlgrey_2.u_pinmux_aon.lc_jtag_i &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.rv_jtag_i    == top_level_upec.top_earlgrey_2.u_pinmux_aon.rv_jtag_i &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dft_jtag_i   == top_level_upec.top_earlgrey_2.u_pinmux_aon.dft_jtag_i    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dft_hold_tap_sel_i   == top_level_upec.top_earlgrey_2.u_pinmux_aon.dft_hold_tap_sel_i    &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.sleep_en_i   == top_level_upec.top_earlgrey_2.u_pinmux_aon.sleep_en_i    &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.strap_en_i   == top_level_upec.top_earlgrey_2.u_pinmux_aon.strap_en_i    &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.usb_out_of_rst_i == top_level_upec.top_earlgrey_2.u_pinmux_aon.usb_out_of_rst_i  &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.usb_aon_wake_en_i    == top_level_upec.top_earlgrey_2.u_pinmux_aon.usb_aon_wake_en_i &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.usb_aon_wake_ack_i   == top_level_upec.top_earlgrey_2.u_pinmux_aon.usb_aon_wake_ack_i    &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.usb_suspend_i    == top_level_upec.top_earlgrey_2.u_pinmux_aon.usb_suspend_i &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.tl_i == top_level_upec.top_earlgrey_2.u_pinmux_aon.tl_i  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.periph_to_mio_i[52]  == top_level_upec.top_earlgrey_2.u_pinmux_aon.periph_to_mio_i[52]   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.periph_to_mio_i[71:68]  == top_level_upec.top_earlgrey_2.u_pinmux_aon.periph_to_mio_i[71:68]   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.periph_to_mio_oe_i[52]   == top_level_upec.top_earlgrey_2.u_pinmux_aon.periph_to_mio_oe_i[52]    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.periph_to_mio_oe_i[71:68]   == top_level_upec.top_earlgrey_2.u_pinmux_aon.periph_to_mio_oe_i[71:68]    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_in_i == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_in_i  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.periph_to_dio_i[23:22]  == top_level_upec.top_earlgrey_2.u_pinmux_aon.periph_to_dio_i[23:22]   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.periph_to_dio_oe_i[23:22]   == top_level_upec.top_earlgrey_2.u_pinmux_aon.periph_to_dio_oe_i[23:22]    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_in_i == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_in_i  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.scanmode_i   == top_level_upec.top_earlgrey_2.u_pinmux_aon.scanmode_i
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.clk_i    == top_level_upec.top_earlgrey_2.u_pinmux_aon.clk_i &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.clk_aon_i    == top_level_upec.top_earlgrey_2.u_pinmux_aon.clk_aon_i &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.rst_ni   == top_level_upec.top_earlgrey_2.u_pinmux_aon.rst_ni    &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.rst_aon_ni   == top_level_upec.top_earlgrey_2.u_pinmux_aon.rst_aon_ni    &&

    );
endfunction

function automatic output_equivalence_peri_devices();
    output_equivalence_peri_devices = (
//        top_level_upec.top_earlgrey_1.u_uart0.cio_tx_o  == top_level_upec.top_earlgrey_2.u_uart0.cio_tx_o   &&   
//        top_level_upec.top_earlgrey_1.u_uart0.cio_tx_en_o   == top_level_upec.top_earlgrey_2.u_uart0.cio_tx_en_o    &&
        top_level_upec.top_earlgrey_1.u_uart0.intr_tx_watermark_o   == top_level_upec.top_earlgrey_2.u_uart0.intr_tx_watermark_o    &&  
        top_level_upec.top_earlgrey_1.u_uart0.intr_rx_watermark_o   == top_level_upec.top_earlgrey_2.u_uart0.intr_rx_watermark_o    &&  
        top_level_upec.top_earlgrey_1.u_uart0.intr_tx_empty_o   == top_level_upec.top_earlgrey_2.u_uart0.intr_tx_empty_o    &&      
        top_level_upec.top_earlgrey_1.u_uart0.intr_rx_overflow_o    == top_level_upec.top_earlgrey_2.u_uart0.intr_rx_overflow_o &&   
        top_level_upec.top_earlgrey_1.u_uart0.intr_rx_frame_err_o   == top_level_upec.top_earlgrey_2.u_uart0.intr_rx_frame_err_o    &&  
        top_level_upec.top_earlgrey_1.u_uart0.intr_rx_break_err_o   == top_level_upec.top_earlgrey_2.u_uart0.intr_rx_break_err_o    &&  
        top_level_upec.top_earlgrey_1.u_uart0.intr_rx_timeout_o == top_level_upec.top_earlgrey_2.u_uart0.intr_rx_timeout_o  &&    
        top_level_upec.top_earlgrey_1.u_uart0.intr_rx_parity_err_o  == top_level_upec.top_earlgrey_2.u_uart0.intr_rx_parity_err_o   && 
//        top_level_upec.top_earlgrey_1.u_uart0.alert_tx_o    == top_level_upec.top_earlgrey_2.u_uart0.alert_tx_o &&
//        top_level_upec.top_earlgrey_1.u_uart0.tl_o  == top_level_upec.top_earlgrey_2.u_uart0.tl_o   &&

//        top_level_upec.top_earlgrey_1.u_uart1.cio_tx_o  == top_level_upec.top_earlgrey_2.u_uart1.cio_tx_o   &&   
//        top_level_upec.top_earlgrey_1.u_uart1.cio_tx_en_o   == top_level_upec.top_earlgrey_2.u_uart1.cio_tx_en_o    &&
        top_level_upec.top_earlgrey_1.u_uart1.intr_tx_watermark_o   == top_level_upec.top_earlgrey_2.u_uart1.intr_tx_watermark_o    &&  
        top_level_upec.top_earlgrey_1.u_uart1.intr_rx_watermark_o   == top_level_upec.top_earlgrey_2.u_uart1.intr_rx_watermark_o    &&  
        top_level_upec.top_earlgrey_1.u_uart1.intr_tx_empty_o   == top_level_upec.top_earlgrey_2.u_uart1.intr_tx_empty_o    &&      
        top_level_upec.top_earlgrey_1.u_uart1.intr_rx_overflow_o    == top_level_upec.top_earlgrey_2.u_uart1.intr_rx_overflow_o &&   
        top_level_upec.top_earlgrey_1.u_uart1.intr_rx_frame_err_o   == top_level_upec.top_earlgrey_2.u_uart1.intr_rx_frame_err_o    &&  
        top_level_upec.top_earlgrey_1.u_uart1.intr_rx_break_err_o   == top_level_upec.top_earlgrey_2.u_uart1.intr_rx_break_err_o    &&  
        top_level_upec.top_earlgrey_1.u_uart1.intr_rx_timeout_o == top_level_upec.top_earlgrey_2.u_uart1.intr_rx_timeout_o  &&    
        top_level_upec.top_earlgrey_1.u_uart1.intr_rx_parity_err_o  == top_level_upec.top_earlgrey_2.u_uart1.intr_rx_parity_err_o   && 
//        top_level_upec.top_earlgrey_1.u_uart1.alert_tx_o    == top_level_upec.top_earlgrey_2.u_uart1.alert_tx_o &&
//        top_level_upec.top_earlgrey_1.u_uart1.tl_o  == top_level_upec.top_earlgrey_2.u_uart1.tl_o   &&

//        top_level_upec.top_earlgrey_1.u_uart2.cio_tx_o  == top_level_upec.top_earlgrey_2.u_uart2.cio_tx_o   &&   
//        top_level_upec.top_earlgrey_1.u_uart2.cio_tx_en_o   == top_level_upec.top_earlgrey_2.u_uart2.cio_tx_en_o    &&
        top_level_upec.top_earlgrey_1.u_uart2.intr_tx_watermark_o   == top_level_upec.top_earlgrey_2.u_uart2.intr_tx_watermark_o    &&  
        top_level_upec.top_earlgrey_1.u_uart2.intr_rx_watermark_o   == top_level_upec.top_earlgrey_2.u_uart2.intr_rx_watermark_o    &&  
        top_level_upec.top_earlgrey_1.u_uart2.intr_tx_empty_o   == top_level_upec.top_earlgrey_2.u_uart2.intr_tx_empty_o    &&      
        top_level_upec.top_earlgrey_1.u_uart2.intr_rx_overflow_o    == top_level_upec.top_earlgrey_2.u_uart2.intr_rx_overflow_o &&   
        top_level_upec.top_earlgrey_1.u_uart2.intr_rx_frame_err_o   == top_level_upec.top_earlgrey_2.u_uart2.intr_rx_frame_err_o    &&  
        top_level_upec.top_earlgrey_1.u_uart2.intr_rx_break_err_o   == top_level_upec.top_earlgrey_2.u_uart2.intr_rx_break_err_o    &&  
        top_level_upec.top_earlgrey_1.u_uart2.intr_rx_timeout_o == top_level_upec.top_earlgrey_2.u_uart2.intr_rx_timeout_o  &&    
        top_level_upec.top_earlgrey_1.u_uart2.intr_rx_parity_err_o  == top_level_upec.top_earlgrey_2.u_uart2.intr_rx_parity_err_o   && 
//        top_level_upec.top_earlgrey_1.u_uart2.alert_tx_o    == top_level_upec.top_earlgrey_2.u_uart2.alert_tx_o &&
//        top_level_upec.top_earlgrey_1.u_uart2.tl_o  == top_level_upec.top_earlgrey_2.u_uart2.tl_o   &&

//        top_level_upec.top_earlgrey_1.u_uart3.cio_tx_o  == top_level_upec.top_earlgrey_2.u_uart3.cio_tx_o   &&   
//        top_level_upec.top_earlgrey_1.u_uart3.cio_tx_en_o   == top_level_upec.top_earlgrey_2.u_uart3.cio_tx_en_o    &&
        top_level_upec.top_earlgrey_1.u_uart3.intr_tx_watermark_o   == top_level_upec.top_earlgrey_2.u_uart3.intr_tx_watermark_o    &&  
        top_level_upec.top_earlgrey_1.u_uart3.intr_rx_watermark_o   == top_level_upec.top_earlgrey_2.u_uart3.intr_rx_watermark_o    &&  
        top_level_upec.top_earlgrey_1.u_uart3.intr_tx_empty_o   == top_level_upec.top_earlgrey_2.u_uart3.intr_tx_empty_o    &&      
        top_level_upec.top_earlgrey_1.u_uart3.intr_rx_overflow_o    == top_level_upec.top_earlgrey_2.u_uart3.intr_rx_overflow_o &&   
        top_level_upec.top_earlgrey_1.u_uart3.intr_rx_frame_err_o   == top_level_upec.top_earlgrey_2.u_uart3.intr_rx_frame_err_o    &&  
        top_level_upec.top_earlgrey_1.u_uart3.intr_rx_break_err_o   == top_level_upec.top_earlgrey_2.u_uart3.intr_rx_break_err_o    &&  
        top_level_upec.top_earlgrey_1.u_uart3.intr_rx_timeout_o == top_level_upec.top_earlgrey_2.u_uart3.intr_rx_timeout_o  &&    
        top_level_upec.top_earlgrey_1.u_uart3.intr_rx_parity_err_o  == top_level_upec.top_earlgrey_2.u_uart3.intr_rx_parity_err_o   && 
//        top_level_upec.top_earlgrey_1.u_uart3.alert_tx_o    == top_level_upec.top_earlgrey_2.u_uart3.alert_tx_o &&
//        top_level_upec.top_earlgrey_1.u_uart3.tl_o  == top_level_upec.top_earlgrey_2.u_uart3.tl_o   &&

//        top_level_upec.top_earlgrey_1.u_spi_host0.cio_sck_o == top_level_upec.top_earlgrey_2.u_spi_host0.cio_sck_o  &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.cio_sck_en_o  == top_level_upec.top_earlgrey_2.u_spi_host0.cio_sck_en_o   &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.cio_csb_o == top_level_upec.top_earlgrey_2.u_spi_host0.cio_csb_o  &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.cio_csb_en_o  == top_level_upec.top_earlgrey_2.u_spi_host0.cio_csb_en_o   &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.cio_sd_o  == top_level_upec.top_earlgrey_2.u_spi_host0.cio_sd_o   &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.cio_sd_en_o   == top_level_upec.top_earlgrey_2.u_spi_host0.cio_sd_en_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.intr_error_o  == top_level_upec.top_earlgrey_2.u_spi_host0.intr_error_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.intr_spi_event_o  == top_level_upec.top_earlgrey_2.u_spi_host0.intr_spi_event_o   &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.alert_tx_o    == top_level_upec.top_earlgrey_2.u_spi_host0.alert_tx_o &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.passthrough_o == top_level_upec.top_earlgrey_2.u_spi_host0.passthrough_o  &&
//        top_level_upec.top_earlgrey_1.u_spi_host0.tl_o  == top_level_upec.top_earlgrey_2.u_spi_host0.tl_o   &&

//        top_level_upec.top_earlgrey_1.u_spi_host1.cio_sck_o == top_level_upec.top_earlgrey_2.u_spi_host1.cio_sck_o  &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.cio_sck_en_o  == top_level_upec.top_earlgrey_2.u_spi_host1.cio_sck_en_o   &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.cio_csb_o == top_level_upec.top_earlgrey_2.u_spi_host1.cio_csb_o  &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.cio_csb_en_o  == top_level_upec.top_earlgrey_2.u_spi_host1.cio_csb_en_o   &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.cio_sd_o  == top_level_upec.top_earlgrey_2.u_spi_host1.cio_sd_o   &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.cio_sd_en_o   == top_level_upec.top_earlgrey_2.u_spi_host1.cio_sd_en_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.intr_error_o  == top_level_upec.top_earlgrey_2.u_spi_host1.intr_error_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.intr_spi_event_o  == top_level_upec.top_earlgrey_2.u_spi_host1.intr_spi_event_o   &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.alert_tx_o    == top_level_upec.top_earlgrey_2.u_spi_host1.alert_tx_o &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.passthrough_o == top_level_upec.top_earlgrey_2.u_spi_host1.passthrough_o  &&
//        top_level_upec.top_earlgrey_1.u_spi_host1.tl_o  == top_level_upec.top_earlgrey_2.u_spi_host1.tl_o   &&
        

//        top_level_upec.top_earlgrey_1.u_spi_device.cio_sd_o == top_level_upec.top_earlgrey_2.u_spi_device.cio_sd_o  &&
//        top_level_upec.top_earlgrey_1.u_spi_device.cio_sd_en_o  == top_level_upec.top_earlgrey_2.u_spi_device.cio_sd_en_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.intr_rxf_o   == top_level_upec.top_earlgrey_2.u_spi_device.intr_rxf_o    &&
        top_level_upec.top_earlgrey_1.u_spi_device.intr_rxlvl_o == top_level_upec.top_earlgrey_2.u_spi_device.intr_rxlvl_o  &&
        top_level_upec.top_earlgrey_1.u_spi_device.intr_txlvl_o == top_level_upec.top_earlgrey_2.u_spi_device.intr_txlvl_o  &&
        top_level_upec.top_earlgrey_1.u_spi_device.intr_rxerr_o == top_level_upec.top_earlgrey_2.u_spi_device.intr_rxerr_o  &&
        top_level_upec.top_earlgrey_1.u_spi_device.intr_rxoverflow_o    == top_level_upec.top_earlgrey_2.u_spi_device.intr_rxoverflow_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.intr_txunderflow_o   == top_level_upec.top_earlgrey_2.u_spi_device.intr_txunderflow_o    &&
//        top_level_upec.top_earlgrey_1.u_spi_device.alert_tx_o   == top_level_upec.top_earlgrey_2.u_spi_device.alert_tx_o    &&
//        top_level_upec.top_earlgrey_1.u_spi_device.passthrough_o    == top_level_upec.top_earlgrey_2.u_spi_device.passthrough_o &&
//        top_level_upec.top_earlgrey_1.u_spi_device.tl_o == top_level_upec.top_earlgrey_2.u_spi_device.tl_o  &&

//        top_level_upec.top_earlgrey_1.u_usbdev.cio_se0_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_se0_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_se0_en_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_se0_en_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_dp_pullup_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_dp_pullup_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_dp_pullup_en_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_dp_pullup_en_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_dn_pullup_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_dn_pullup_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_dn_pullup_en_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_dn_pullup_en_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_tx_mode_se_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_tx_mode_se_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_tx_mode_se_en_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_tx_mode_se_en_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_suspend_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_suspend_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_suspend_en_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_suspend_en_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_rx_enable_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_rx_enable_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_rx_enable_en_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_rx_enable_en_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_d_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_d_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_d_en_o   == top_level_upec.top_earlgrey_2.u_usbdev.cio_d_en_o    &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_dp_o == top_level_upec.top_earlgrey_2.u_usbdev.cio_dp_o  &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_dp_en_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_dp_en_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_dn_o == top_level_upec.top_earlgrey_2.u_usbdev.cio_dn_o  &&
//        top_level_upec.top_earlgrey_1.u_usbdev.cio_dn_en_o  == top_level_upec.top_earlgrey_2.u_usbdev.cio_dn_en_o   && 
        top_level_upec.top_earlgrey_1.u_usbdev.intr_pkt_received_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_pkt_received_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_pkt_sent_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_pkt_sent_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_disconnected_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_disconnected_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_host_lost_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_host_lost_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_reset_o    == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_reset_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_suspend_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_suspend_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_resume_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_resume_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_av_empty_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_av_empty_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_full_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_full_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_av_overflow_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_av_overflow_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_in_err_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_in_err_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_crc_err_o    == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_crc_err_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_pid_err_o    == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_pid_err_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_bitstuff_err_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_bitstuff_err_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_frame_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_frame_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_connected_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_connected_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_out_err_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_out_err_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usb_ref_val_o    == top_level_upec.top_earlgrey_2.u_usbdev.usb_ref_val_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usb_ref_pulse_o  == top_level_upec.top_earlgrey_2.u_usbdev.usb_ref_pulse_o   &&
//        top_level_upec.top_earlgrey_1.u_usbdev.usb_out_of_rst_o == top_level_upec.top_earlgrey_2.u_usbdev.usb_out_of_rst_o  &&
//        top_level_upec.top_earlgrey_1.u_usbdev.usb_aon_wake_en_o    == top_level_upec.top_earlgrey_2.u_usbdev.usb_aon_wake_en_o &&
//        top_level_upec.top_earlgrey_1.u_usbdev.usb_aon_wake_ack_o   == top_level_upec.top_earlgrey_2.u_usbdev.usb_aon_wake_ack_o    &&
//        top_level_upec.top_earlgrey_1.u_usbdev.usb_suspend_o    == top_level_upec.top_earlgrey_2.u_usbdev.usb_suspend_o &&
//        top_level_upec.top_earlgrey_1.u_usbdev.tl_o    == top_level_upec.top_earlgrey_2.u_usbdev.tl_o &&

//        top_level_upec.top_earlgrey_1.u_gpio.cio_gpio_o == top_level_upec.top_earlgrey_2.u_gpio.cio_gpio_o  &&
//        top_level_upec.top_earlgrey_1.u_gpio.cio_gpio_en_o  == top_level_upec.top_earlgrey_2.u_gpio.cio_gpio_en_o   &&
        top_level_upec.top_earlgrey_1.u_gpio.intr_gpio_o    == top_level_upec.top_earlgrey_2.u_gpio.intr_gpio_o &&
//        top_level_upec.top_earlgrey_1.u_gpio.alert_tx_o == top_level_upec.top_earlgrey_2.u_gpio.alert_tx_o  &&
//        top_level_upec.top_earlgrey_1.u_gpio.tl_o   == top_level_upec.top_earlgrey_2.u_gpio.tl_o    &&

//        top_level_upec.top_earlgrey_1.u_i2c0.cio_sda_o  == top_level_upec.top_earlgrey_2.u_i2c0.cio_sda_o   &&
//        top_level_upec.top_earlgrey_1.u_i2c0.cio_sda_en_o   == top_level_upec.top_earlgrey_2.u_i2c0.cio_sda_en_o    &&
//        top_level_upec.top_earlgrey_1.u_i2c0.cio_scl_o  == top_level_upec.top_earlgrey_2.u_i2c0.cio_scl_o   &&
//        top_level_upec.top_earlgrey_1.u_i2c0.cio_scl_en_o   == top_level_upec.top_earlgrey_2.u_i2c0.cio_scl_en_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_fmt_watermark_o   == top_level_upec.top_earlgrey_2.u_i2c0.intr_fmt_watermark_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_rx_watermark_o    == top_level_upec.top_earlgrey_2.u_i2c0.intr_rx_watermark_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_fmt_overflow_o    == top_level_upec.top_earlgrey_2.u_i2c0.intr_fmt_overflow_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_rx_overflow_o == top_level_upec.top_earlgrey_2.u_i2c0.intr_rx_overflow_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_nak_o == top_level_upec.top_earlgrey_2.u_i2c0.intr_nak_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_scl_interference_o    == top_level_upec.top_earlgrey_2.u_i2c0.intr_scl_interference_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_sda_interference_o    == top_level_upec.top_earlgrey_2.u_i2c0.intr_sda_interference_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_stretch_timeout_o == top_level_upec.top_earlgrey_2.u_i2c0.intr_stretch_timeout_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_sda_unstable_o    == top_level_upec.top_earlgrey_2.u_i2c0.intr_sda_unstable_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_trans_complete_o  == top_level_upec.top_earlgrey_2.u_i2c0.intr_trans_complete_o   &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_tx_empty_o    == top_level_upec.top_earlgrey_2.u_i2c0.intr_tx_empty_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_tx_nonempty_o == top_level_upec.top_earlgrey_2.u_i2c0.intr_tx_nonempty_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_tx_overflow_o == top_level_upec.top_earlgrey_2.u_i2c0.intr_tx_overflow_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_acq_overflow_o    == top_level_upec.top_earlgrey_2.u_i2c0.intr_acq_overflow_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_ack_stop_o    == top_level_upec.top_earlgrey_2.u_i2c0.intr_ack_stop_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.intr_host_timeout_o    == top_level_upec.top_earlgrey_2.u_i2c0.intr_host_timeout_o &&
//        top_level_upec.top_earlgrey_1.u_i2c0.alert_tx_o == top_level_upec.top_earlgrey_2.u_i2c0.alert_tx_o  &&
//        top_level_upec.top_earlgrey_1.u_i2c0.tl_o   == top_level_upec.top_earlgrey_2.u_i2c0.tl_o    &&

//        top_level_upec.top_earlgrey_1.u_i2c1.cio_sda_o  == top_level_upec.top_earlgrey_2.u_i2c1.cio_sda_o   &&
//        top_level_upec.top_earlgrey_1.u_i2c1.cio_sda_en_o   == top_level_upec.top_earlgrey_2.u_i2c1.cio_sda_en_o    &&
//        top_level_upec.top_earlgrey_1.u_i2c1.cio_scl_o  == top_level_upec.top_earlgrey_2.u_i2c1.cio_scl_o   &&
//        top_level_upec.top_earlgrey_1.u_i2c1.cio_scl_en_o   == top_level_upec.top_earlgrey_2.u_i2c1.cio_scl_en_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_fmt_watermark_o   == top_level_upec.top_earlgrey_2.u_i2c1.intr_fmt_watermark_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_rx_watermark_o    == top_level_upec.top_earlgrey_2.u_i2c1.intr_rx_watermark_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_fmt_overflow_o    == top_level_upec.top_earlgrey_2.u_i2c1.intr_fmt_overflow_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_rx_overflow_o == top_level_upec.top_earlgrey_2.u_i2c1.intr_rx_overflow_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_nak_o == top_level_upec.top_earlgrey_2.u_i2c1.intr_nak_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_scl_interference_o    == top_level_upec.top_earlgrey_2.u_i2c1.intr_scl_interference_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_sda_interference_o    == top_level_upec.top_earlgrey_2.u_i2c1.intr_sda_interference_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_stretch_timeout_o == top_level_upec.top_earlgrey_2.u_i2c1.intr_stretch_timeout_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_sda_unstable_o    == top_level_upec.top_earlgrey_2.u_i2c1.intr_sda_unstable_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_trans_complete_o  == top_level_upec.top_earlgrey_2.u_i2c1.intr_trans_complete_o   &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_tx_empty_o    == top_level_upec.top_earlgrey_2.u_i2c1.intr_tx_empty_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_tx_nonempty_o == top_level_upec.top_earlgrey_2.u_i2c1.intr_tx_nonempty_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_tx_overflow_o == top_level_upec.top_earlgrey_2.u_i2c1.intr_tx_overflow_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_acq_overflow_o    == top_level_upec.top_earlgrey_2.u_i2c1.intr_acq_overflow_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_ack_stop_o    == top_level_upec.top_earlgrey_2.u_i2c1.intr_ack_stop_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.intr_host_timeout_o    == top_level_upec.top_earlgrey_2.u_i2c1.intr_host_timeout_o &&
//        top_level_upec.top_earlgrey_1.u_i2c1.alert_tx_o == top_level_upec.top_earlgrey_2.u_i2c1.alert_tx_o  &&
//        top_level_upec.top_earlgrey_1.u_i2c1.tl_o   == top_level_upec.top_earlgrey_2.u_i2c1.tl_o    &&

//        top_level_upec.top_earlgrey_1.u_i2c2.cio_sda_o  == top_level_upec.top_earlgrey_2.u_i2c2.cio_sda_o   &&
//        top_level_upec.top_earlgrey_1.u_i2c2.cio_sda_en_o   == top_level_upec.top_earlgrey_2.u_i2c2.cio_sda_en_o    &&
//        top_level_upec.top_earlgrey_1.u_i2c2.cio_scl_o  == top_level_upec.top_earlgrey_2.u_i2c2.cio_scl_o   &&
//        top_level_upec.top_earlgrey_1.u_i2c2.cio_scl_en_o   == top_level_upec.top_earlgrey_2.u_i2c2.cio_scl_en_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_fmt_watermark_o   == top_level_upec.top_earlgrey_2.u_i2c2.intr_fmt_watermark_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_rx_watermark_o    == top_level_upec.top_earlgrey_2.u_i2c2.intr_rx_watermark_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_fmt_overflow_o    == top_level_upec.top_earlgrey_2.u_i2c2.intr_fmt_overflow_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_rx_overflow_o == top_level_upec.top_earlgrey_2.u_i2c2.intr_rx_overflow_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_nak_o == top_level_upec.top_earlgrey_2.u_i2c2.intr_nak_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_scl_interference_o    == top_level_upec.top_earlgrey_2.u_i2c2.intr_scl_interference_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_sda_interference_o    == top_level_upec.top_earlgrey_2.u_i2c2.intr_sda_interference_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_stretch_timeout_o == top_level_upec.top_earlgrey_2.u_i2c2.intr_stretch_timeout_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_sda_unstable_o    == top_level_upec.top_earlgrey_2.u_i2c2.intr_sda_unstable_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_trans_complete_o  == top_level_upec.top_earlgrey_2.u_i2c2.intr_trans_complete_o   &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_tx_empty_o    == top_level_upec.top_earlgrey_2.u_i2c2.intr_tx_empty_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_tx_nonempty_o == top_level_upec.top_earlgrey_2.u_i2c2.intr_tx_nonempty_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_tx_overflow_o == top_level_upec.top_earlgrey_2.u_i2c2.intr_tx_overflow_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_acq_overflow_o    == top_level_upec.top_earlgrey_2.u_i2c2.intr_acq_overflow_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_ack_stop_o    == top_level_upec.top_earlgrey_2.u_i2c2.intr_ack_stop_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.intr_host_timeout_o    == top_level_upec.top_earlgrey_2.u_i2c2.intr_host_timeout_o &&
//        top_level_upec.top_earlgrey_1.u_i2c2.alert_tx_o == top_level_upec.top_earlgrey_2.u_i2c2.alert_tx_o  &&
//        top_level_upec.top_earlgrey_1.u_i2c2.tl_o   == top_level_upec.top_earlgrey_2.u_i2c2.tl_o    &&

//        top_level_upec.top_earlgrey_1.u_pwm_aon.cio_pwm_o   == top_level_upec.top_earlgrey_2.u_pwm_aon.cio_pwm_o    &&
//        top_level_upec.top_earlgrey_1.u_pwm_aon.cio_pwm_en_o    == top_level_upec.top_earlgrey_2.u_pwm_aon.cio_pwm_en_o &&
//        top_level_upec.top_earlgrey_1.u_pwm_aon.tl_o    == top_level_upec.top_earlgrey_2.u_pwm_aon.tl_o &&

        top_level_upec.top_earlgrey_1.u_clkmgr_aon.clocks_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.clocks_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.ast_clk_byp_req_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.ast_clk_byp_req_o &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.lc_clk_byp_ack_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.lc_clk_byp_ack_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.jitter_en_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.jitter_en_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.clocks_ast_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.clocks_ast_o  &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.pwr_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.pwr_o &&
//        top_level_upec.top_earlgrey_1.u_clkmgr_aon.tl_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.tl_o  &&

        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.intr_wakeup_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.intr_wakeup_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_ast_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_ast_o &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_rst_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_rst_o &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_clk_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_clk_o &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_otp_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_otp_o &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.pwr_lc_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.pwr_lc_o  &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.esc_rst_rx_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.esc_rst_rx_o  &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.strap_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.strap_o   &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.low_power_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.low_power_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.fetch_en_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.fetch_en_o    &&
//        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.tl_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.tl_o  &&

        top_level_upec.top_earlgrey_1.u_rv_timer.intr_timer_expired_0_0_o   == top_level_upec.top_earlgrey_2.u_rv_timer.intr_timer_expired_0_0_o    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.intr_timer_expired_1_0_o   == top_level_upec.top_earlgrey_2.u_rv_timer.intr_timer_expired_1_0_o    &&
//        top_level_upec.top_earlgrey_1.u_rv_timer.tl_o   == top_level_upec.top_earlgrey_2.u_rv_timer.tl_o    &&

        top_level_upec.top_earlgrey_1.u_alert_handler.intr_classa_o == top_level_upec.top_earlgrey_2.u_alert_handler.intr_classa_o  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.intr_classb_o == top_level_upec.top_earlgrey_2.u_alert_handler.intr_classb_o  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.intr_classc_o == top_level_upec.top_earlgrey_2.u_alert_handler.intr_classc_o  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.intr_classd_o == top_level_upec.top_earlgrey_2.u_alert_handler.intr_classd_o  &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.crashdump_o   == top_level_upec.top_earlgrey_2.u_alert_handler.crashdump_o    &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.edn_o == top_level_upec.top_earlgrey_2.u_alert_handler.edn_o  &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.esc_tx_o  == top_level_upec.top_earlgrey_2.u_alert_handler.esc_tx_o   &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.tl_o  == top_level_upec.top_earlgrey_2.u_alert_handler.tl_o   &&
//        top_level_upec.top_earlgrey_1.u_alert_handler.alert_rx_o[31:0]    == top_level_upec.top_earlgrey_2.u_alert_handler.alert_rx_o[31:0] &&
        top_level_upec.top_earlgrey_1.u_alert_handler.alert_rx_o[51:32]    == top_level_upec.top_earlgrey_2.u_alert_handler.alert_rx_o[51:32]   &&

        top_level_upec.top_earlgrey_1.u_aon_timer_aon.intr_wkup_timer_expired_o == top_level_upec.top_earlgrey_2.u_aon_timer_aon.intr_wkup_timer_expired_o  &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.intr_wdog_timer_bark_o    == top_level_upec.top_earlgrey_2.u_aon_timer_aon.intr_wdog_timer_bark_o &&
//        top_level_upec.top_earlgrey_1.u_aon_timer_aon.aon_timer_wkup_req_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.aon_timer_wkup_req_o   &&
//        top_level_upec.top_earlgrey_1.u_aon_timer_aon.aon_timer_rst_req_o   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.aon_timer_rst_req_o    &&
//        top_level_upec.top_earlgrey_1.u_aon_timer_aon.tl_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.tl_o   &&

        top_level_upec.top_earlgrey_1.u_otp_ctrl.intr_otp_operation_done_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.intr_otp_operation_done_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.intr_otp_error_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.intr_otp_error_o    &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.alert_tx_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.alert_tx_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.otp_ast_pwr_seq_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.otp_ast_pwr_seq_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.otp_alert_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.otp_alert_o &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.edn_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.edn_o   &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.pwr_otp_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.pwr_otp_o   &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.lc_otp_program_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.lc_otp_program_o    &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.otp_lc_data_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.otp_lc_data_o   &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.otp_keymgr_key_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.otp_keymgr_key_o    &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.flash_otp_key_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.flash_otp_key_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.sram_otp_key_o[0] == top_level_upec.top_earlgrey_2.u_otp_ctrl.sram_otp_key_o[0]  &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.sram_otp_key_o[1] == top_level_upec.top_earlgrey_2.u_otp_ctrl.sram_otp_key_o[1]  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.otbn_otp_key_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.otbn_otp_key_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.otp_hw_cfg_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.otp_hw_cfg_o    &&
//        top_level_upec.top_earlgrey_1.u_otp_ctrl.tl_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.tl_o    &&

//        top_level_upec.top_earlgrey_1.u_lc_ctrl.alert_tx_o    == top_level_upec.top_earlgrey_2.lc_ctrl.alert_tx_o &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.jtag_o    == top_level_upec.top_earlgrey_2.lc_ctrl.jtag_o &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.esc_wipe_secrets_rx_o == top_level_upec.top_earlgrey_2.lc_ctrl.esc_wipe_secrets_rx_o  &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.esc_scrap_state_rx_o  == top_level_upec.top_earlgrey_2.lc_ctrl.esc_scrap_state_rx_o   &&
 //       top_level_upec.top_earlgrey_1.u_lc_ctrl.pwr_lc_o  == top_level_upec.top_earlgrey_2.lc_ctrl.pwr_lc_o   &&
  //      top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_otp_program_o  == top_level_upec.top_earlgrey_2.lc_ctrl.lc_otp_program_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.kmac_data_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.kmac_data_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_dft_en_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_dft_en_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_nvm_debug_en_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_nvm_debug_en_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_hw_debug_en_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_hw_debug_en_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_cpu_en_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_cpu_en_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_keymgr_en_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_keymgr_en_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_escalate_en_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_escalate_en_o   &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_clk_byp_req_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_clk_byp_req_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_flash_rma_req_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_flash_rma_req_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_flash_rma_seed_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_flash_rma_seed_o    &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_check_byp_en_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_check_byp_en_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_creator_seed_sw_rw_en_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_creator_seed_sw_rw_en_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_owner_seed_sw_rw_en_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_owner_seed_sw_rw_en_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_iso_part_sw_rd_en_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_iso_part_sw_rd_en_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_iso_part_sw_wr_en_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_iso_part_sw_wr_en_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_seed_hw_rd_en_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_seed_hw_rd_en_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_keymgr_div_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_keymgr_div_o    &&
//        top_level_upec.top_earlgrey_1.u_lc_ctrl.tl_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.tl_o   &&

//        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.tl_o == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.tl_o  &&
////        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.req_o    == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.req_o &&
////        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.req_type_o   == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.req_type_o    &&
////        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.we_o == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.we_o  &&
////        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.addr_o   == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.addr_o    &&
////        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.wdata_o  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.wdata_o   &&
////        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.wmask_o  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.wmask_o   &&
////        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.intg_error_o == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.intg_error_o  &&

//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.alert_tx_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.alert_tx_o &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.sram_otp_key_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.sram_otp_key_o &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.sram_scr_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.sram_scr_o &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.sram_scr_init_o   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.sram_scr_init_o    &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.en_ifetch_o   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.en_ifetch_o    &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.tl_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.tl_o   &&

//        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.cio_ast_debug_out_o == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.cio_ast_debug_out_o  &&
//        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.cio_ast_debug_out_en_o  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.cio_ast_debug_out_en_o   &&
//        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.alert_tx_o  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.alert_tx_o   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.ast_alert_o == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.ast_alert_o  &&
//        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.tl_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.tl_o &&

//        top_level_upec.top_earlgrey_1.u_pattgen.cio_pda0_tx_o   == top_level_upec.top_earlgrey_2.u_pattgen.cio_pda0_tx_o    &&
//        top_level_upec.top_earlgrey_1.u_pattgen.cio_pda0_tx_en_o    == top_level_upec.top_earlgrey_2.u_pattgen.cio_pda0_tx_en_o &&
//        top_level_upec.top_earlgrey_1.u_pattgen.cio_pcl0_tx_o   == top_level_upec.top_earlgrey_2.u_pattgen.cio_pcl0_tx_o    &&
//        top_level_upec.top_earlgrey_1.u_pattgen.cio_pcl0_tx_en_o    == top_level_upec.top_earlgrey_2.u_pattgen.cio_pcl0_tx_en_o &&
//        top_level_upec.top_earlgrey_1.u_pattgen.cio_pda1_tx_o   == top_level_upec.top_earlgrey_2.u_pattgen.cio_pda1_tx_o    &&
//        top_level_upec.top_earlgrey_1.u_pattgen.cio_pda1_tx_en_o    == top_level_upec.top_earlgrey_2.u_pattgen.cio_pda1_tx_en_o &&
//        top_level_upec.top_earlgrey_1.u_pattgen.cio_pcl1_tx_o   == top_level_upec.top_earlgrey_2.u_pattgen.cio_pcl1_tx_o    &&
//        top_level_upec.top_earlgrey_1.u_pattgen.cio_pcl1_tx_en_o    == top_level_upec.top_earlgrey_2.u_pattgen.cio_pcl1_tx_en_o &&
        top_level_upec.top_earlgrey_1.u_pattgen.intr_done_ch0_o == top_level_upec.top_earlgrey_2.u_pattgen.intr_done_ch0_o  &&
        top_level_upec.top_earlgrey_1.u_pattgen.intr_done_ch1_o == top_level_upec.top_earlgrey_2.u_pattgen.intr_done_ch1_o  &&
//        top_level_upec.top_earlgrey_1.u_pattgen.alert_tx_o  == top_level_upec.top_earlgrey_2.u_pattgen.alert_tx_o   &&
//        top_level_upec.top_earlgrey_1.u_pattgen.tl_o    == top_level_upec.top_earlgrey_2.u_pattgen.tl_o &&

//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_bat_disable_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_bat_disable_o    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_bat_disable_en_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_bat_disable_en_o &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_ec_rst_out_l_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_ec_rst_out_l_o   &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_ec_rst_out_l_en_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_ec_rst_out_l_en_o    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_key0_out_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_key0_out_o   &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_key0_out_en_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_key0_out_en_o    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_key1_out_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_key1_out_o   &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_key1_out_en_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_key1_out_en_o    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_key2_out_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_key2_out_o   &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_key2_out_en_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_key2_out_en_o    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_pwrb_out_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_pwrb_out_o   &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.cio_pwrb_out_en_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.cio_pwrb_out_en_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.intr_sysrst_ctrl_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.intr_sysrst_ctrl_o   &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.gsc_wk_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.gsc_wk_o &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.gsc_rst_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.gsc_rst_o    &&
//        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.tl_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.tl_o &&

//        top_level_upec.top_earlgrey_1.u_pinmux_aon.alert_tx_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.alert_tx_o    &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.lc_jtag_o    == top_level_upec.top_earlgrey_2.u_pinmux_aon.lc_jtag_o &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.rv_jtag_o    == top_level_upec.top_earlgrey_2.u_pinmux_aon.rv_jtag_o &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dft_jtag_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.dft_jtag_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dft_strap_test_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.dft_strap_test_o  &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.aon_wkup_req_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.aon_wkup_req_o    &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.usb_wkup_req_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.usb_wkup_req_o    &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.usb_state_debug_o    == top_level_upec.top_earlgrey_2.u_pinmux_aon.usb_state_debug_o &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.tl_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.tl_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_to_periph_o[54:46]  == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_to_periph_o[54:46]   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_attr_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_attr_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_out_o    == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_out_o &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_oe_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_oe_o  &&
//        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_to_periph_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_to_periph_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_attr_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_attr_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_out_o    == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_out_o &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_oe_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_oe_o
    );
endfunction

function automatic micro_soc_state_equivalence_peri_devices();
    micro_soc_state_equivalence_peri_devices = (
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn0_max_v == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn0_max_v  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn0_min_v == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn0_min_v  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn1_max_v == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn1_max_v  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn1_min_v == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn1_min_v  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_lp_sample_cnt  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_lp_sample_cnt   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_np_sample_cnt  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_np_sample_cnt   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_pwrup_time == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_pwrup_time  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_wakeup_time    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_wakeup_time &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.dst_level_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.src_level  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.src_level   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.adc_ctrl_match_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.adc_ctrl_match_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn0_val    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn0_val &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn0_val_we == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn0_val_we  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn1_val    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn1_val &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn1_val_we == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn1_val_we  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.fsm_state_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.fsm_state_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.lp_sample_cnt_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.lp_sample_cnt_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.np_sample_cnt_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.np_sample_cnt_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.pwrup_timer_cnt_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.pwrup_timer_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.trigger_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.trigger_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.wakeup_timer_cnt_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.wakeup_timer_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_adc_ctrl_intr_o.intr_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_adc_ctrl_intr_o.intr_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.dst_level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.src_level    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.src_level &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.dst_level_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.src_level == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.src_level  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.dst_level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.src_level    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.src_level &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.dst_level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.src_level    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.src_level &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.dst_level_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.src_level  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.src_level   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.dst_level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.src_level    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.src_level &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.dst_level_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.src_level == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.src_level  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.dst_level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.src_level    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.src_level &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_adc_enable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_adc_enable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_adc_enable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_adc_enable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.storage == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.storage  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.storage == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.storage  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_fsm_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_fsm_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_fsm_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_fsm_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en3.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en3.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en3.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en3.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en5.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en5.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en5.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en5.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en6.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en6.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en6.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en6.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en7.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en7.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en7.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en7.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_intr_en.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_intr_en.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_intr_en.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_intr_en.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_gray_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_sync_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_sync_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_wptr_gray_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_wptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_wptr_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_wptr_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.storage   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.storage    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en3.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en3.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en3.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en3.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en5.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en5.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en5.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en5.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en6.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en6.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en6.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en6.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en7.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en7.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en7.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en7.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_gray_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_sync_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_sync_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_wptr_gray_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_wptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_wptr_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_wptr_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.storage  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.storage   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.dst_level_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.src_level   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.src_level    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_cond_0.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_cond_0.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_cond_0.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_cond_0.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_max_v_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_max_v_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_max_v_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_max_v_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_min_v_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_min_v_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_min_v_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_min_v_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_cond_1.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_cond_1.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_cond_1.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_cond_1.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_max_v_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_max_v_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_max_v_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_max_v_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_min_v_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_min_v_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_min_v_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_min_v_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_cond_2.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_cond_2.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_cond_2.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_cond_2.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_max_v_2.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_max_v_2.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_max_v_2.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_max_v_2.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_min_v_2.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_min_v_2.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_min_v_2.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_min_v_2.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_cond_3.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_cond_3.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_cond_3.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_cond_3.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_max_v_3.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_max_v_3.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_max_v_3.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_max_v_3.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_min_v_3.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_min_v_3.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_min_v_3.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_min_v_3.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_cond_4.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_cond_4.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_cond_4.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_cond_4.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_max_v_4.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_max_v_4.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_max_v_4.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_max_v_4.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_min_v_4.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_min_v_4.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_min_v_4.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_min_v_4.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_cond_5.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_cond_5.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_cond_5.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_cond_5.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_max_v_5.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_max_v_5.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_max_v_5.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_max_v_5.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_min_v_5.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_min_v_5.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_min_v_5.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_min_v_5.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_cond_6.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_cond_6.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_cond_6.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_cond_6.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_max_v_6.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_max_v_6.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_max_v_6.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_max_v_6.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_min_v_6.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_min_v_6.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_min_v_6.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_min_v_6.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_cond_7.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_cond_7.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_cond_7.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_cond_7.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_max_v_7.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_max_v_7.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_max_v_7.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_max_v_7.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_min_v_7.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_min_v_7.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_min_v_7.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_min_v_7.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_cond_0.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_cond_0.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_cond_0.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_cond_0.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_max_v_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_max_v_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_max_v_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_max_v_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_min_v_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_min_v_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_min_v_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_min_v_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_cond_1.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_cond_1.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_cond_1.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_cond_1.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_max_v_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_max_v_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_max_v_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_max_v_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_min_v_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_min_v_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_min_v_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_min_v_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_cond_2.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_cond_2.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_cond_2.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_cond_2.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_max_v_2.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_max_v_2.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_max_v_2.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_max_v_2.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_min_v_2.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_min_v_2.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_min_v_2.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_min_v_2.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_cond_3.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_cond_3.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_cond_3.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_cond_3.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_max_v_3.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_max_v_3.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_max_v_3.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_max_v_3.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_min_v_3.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_min_v_3.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_min_v_3.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_min_v_3.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_cond_4.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_cond_4.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_cond_4.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_cond_4.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_max_v_4.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_max_v_4.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_max_v_4.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_max_v_4.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_min_v_4.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_min_v_4.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_min_v_4.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_min_v_4.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_cond_5.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_cond_5.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_cond_5.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_cond_5.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_max_v_5.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_max_v_5.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_max_v_5.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_max_v_5.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_min_v_5.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_min_v_5.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_min_v_5.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_min_v_5.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_cond_6.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_cond_6.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_cond_6.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_cond_6.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_max_v_6.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_max_v_6.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_max_v_6.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_max_v_6.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_min_v_6.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_min_v_6.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_min_v_6.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_min_v_6.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_cond_7.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_cond_7.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_cond_7.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_cond_7.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_max_v_7.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_max_v_7.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_max_v_7.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_max_v_7.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_min_v_7.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_min_v_7.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_min_v_7.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_min_v_7.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_ext_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_ext_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_ext_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_ext_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_0.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_0.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_0.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_0.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_ext_0.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_ext_0.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_ext_0.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_ext_0.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_ext_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_ext_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_ext_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_ext_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_1.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_1.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_1.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_1.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_ext_1.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_ext_1.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_ext_1.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_ext_1.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_adc_enable.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_adc_enable.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_adc_enable.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_adc_enable.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_oneshot_mode.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_oneshot_mode.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_oneshot_mode.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_oneshot_mode.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_fsm_rst.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_fsm_rst.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_fsm_rst.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_fsm_rst.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter0_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter0_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter0_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter0_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter1_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter1_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter1_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter1_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter2_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter2_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter2_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter2_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter3_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter3_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter3_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter3_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter4_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter4_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter4_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter4_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter5_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter5_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter5_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter5_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter6_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter6_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter6_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter6_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter7_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter7_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter7_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter7_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_oneshot_intr_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_oneshot_intr_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_oneshot_intr_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_oneshot_intr_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_sink_det.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_sink_det.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_sink_det.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_sink_det.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det_flip.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det_flip.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det_flip.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det_flip.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_3a0_sink_det.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_3a0_sink_det.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_3a0_sink_det.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_3a0_sink_det.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_discon.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_discon.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_discon.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_discon.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_sink_det.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_sink_det.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_sink_det.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_sink_det.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det_flip.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det_flip.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det_flip.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det_flip.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_oneshot.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_oneshot.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_oneshot.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_oneshot.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_lp_sample_ctl.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_lp_sample_ctl.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_lp_sample_ctl.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_lp_sample_ctl.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_lp_mode.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_lp_mode.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_lp_mode.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_lp_mode.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_pwrup_time.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_pwrup_time.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_pwrup_time.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_pwrup_time.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_wakeup_time.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_wakeup_time.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_wakeup_time.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_wakeup_time.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_sample_ctl.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_sample_ctl.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_sample_ctl.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_sample_ctl.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter0_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter0_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter0_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter0_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter1_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter1_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter1_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter1_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter2_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter2_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter2_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter2_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter3_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter3_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter3_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter3_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter4_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter4_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter4_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter4_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter5_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter5_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter5_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter5_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter6_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter6_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter6_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter6_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter7_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter7_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter7_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter7_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_sink_det.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_sink_det.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_sink_det.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_sink_det.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det_flip.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det_flip.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det_flip.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det_flip.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_3a0_sink_det.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_3a0_sink_det.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_3a0_sink_det.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_3a0_sink_det.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_discon.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_discon.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_discon.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_discon.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_sink_det.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_sink_det.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_sink_det.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_sink_det.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det_flip.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det_flip.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det_flip.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det_flip.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_intr_enable.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_intr_enable.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_intr_enable.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_intr_enable.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_intr_state.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_intr_state.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_intr_state.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_intr_state.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[0].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[0].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[0].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[0].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[0].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[0].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[0].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[0].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[0].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[0].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[1].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[1].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[1].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[1].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[1].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[1].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[1].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[1].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[1].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[1].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[2].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[2].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[2].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[2].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[2].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[2].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[2].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[2].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[2].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[2].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[3].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[3].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[3].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[3].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[3].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[3].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[3].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[3].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[3].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[3].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.esc_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.esc_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.esc_req_q1    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.esc_req_q1 &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.u_decode_resp.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.u_decode_resp.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.u_decode_resp.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.u_decode_resp.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.esc_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.esc_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.esc_req_q1    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.esc_req_q1 &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.u_decode_resp.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.u_decode_resp.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.u_decode_resp.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.u_decode_resp.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.esc_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.esc_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.esc_req_q1    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.esc_req_q1 &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.u_decode_resp.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.u_decode_resp.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.u_decode_resp.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.u_decode_resp.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.esc_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.esc_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.esc_req_q1    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.esc_req_q1 &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.u_decode_resp.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.u_decode_resp.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.u_decode_resp.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.u_decode_resp.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.fips_q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.fips_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_packer_fifo.clr_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_packer_fifo.clr_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_packer_fifo.data_q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_packer_fifo.data_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_packer_fifo.depth_q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_packer_fifo.depth_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_packer_fifo.gen_unpack_mode.ptr_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_packer_fifo.gen_unpack_mode.ptr_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs   == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs   == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_cnt[0].u_prim_flop_en.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_cnt[0].u_prim_flop_en.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_cnt[1].u_prim_flop_en.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_cnt[1].u_prim_flop_en.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.cnt_q == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.perturbed_q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.perturbed_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.lfsr_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.lfsr_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.cnt_q == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.perturbed_q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.perturbed_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.lfsr_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.lfsr_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.i_irq_classa.intr_o    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.i_irq_classa.intr_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.i_irq_classb.intr_o    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.i_irq_classb.intr_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.i_irq_classc.intr_o    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.i_irq_classc.intr_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.i_irq_classd.intr_o    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.i_irq_classd.intr_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_10.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_10.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_10.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_10.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_11.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_11.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_11.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_11.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_12.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_12.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_12.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_12.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_13.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_13.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_13.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_13.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_14.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_14.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_14.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_14.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_15.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_15.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_15.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_15.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_16.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_16.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_16.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_16.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_17.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_17.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_17.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_17.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_18.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_18.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_18.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_18.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_19.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_19.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_19.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_19.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_20.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_20.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_20.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_20.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_21.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_21.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_21.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_21.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_22.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_22.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_22.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_22.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_23.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_23.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_23.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_23.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_24.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_24.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_24.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_24.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_25.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_25.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_25.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_25.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_26.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_26.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_26.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_26.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_27.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_27.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_27.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_27.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_28.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_28.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_28.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_28.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_29.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_29.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_29.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_29.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_30.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_30.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_30.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_30.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_31.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_31.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_31.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_31.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_32.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_32.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_32.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_32.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_33.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_33.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_33.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_33.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_34.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_34.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_34.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_34.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_35.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_35.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_35.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_35.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_36.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_36.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_36.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_36.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_37.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_37.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_37.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_37.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_38.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_38.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_38.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_38.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_39.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_39.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_39.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_39.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_4.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_4.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_4.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_4.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_40.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_40.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_40.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_40.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_41.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_41.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_41.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_41.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_42.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_42.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_42.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_42.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_43.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_43.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_43.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_43.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_44.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_44.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_44.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_44.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_45.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_45.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_45.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_45.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_46.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_46.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_46.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_46.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_47.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_47.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_47.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_47.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_48.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_48.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_48.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_48.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_49.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_49.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_49.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_49.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_5.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_5.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_5.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_5.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_50.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_50.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_50.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_50.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_51.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_51.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_51.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_51.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_6.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_6.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_6.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_6.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_7.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_7.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_7.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_7.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_8.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_8.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_8.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_8.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_9.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_9.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_9.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_9.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_10.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_10.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_10.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_10.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_11.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_11.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_11.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_11.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_12.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_12.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_12.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_12.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_13.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_13.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_13.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_13.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_14.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_14.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_14.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_14.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_15.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_15.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_15.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_15.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_16.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_16.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_16.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_16.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_17.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_17.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_17.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_17.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_18.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_18.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_18.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_18.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_19.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_19.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_19.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_19.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_20.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_20.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_20.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_20.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_21.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_21.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_21.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_21.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_22.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_22.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_22.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_22.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_23.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_23.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_23.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_23.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_24.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_24.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_24.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_24.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_25.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_25.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_25.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_25.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_26.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_26.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_26.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_26.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_27.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_27.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_27.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_27.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_28.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_28.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_28.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_28.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_29.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_29.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_29.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_29.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_30.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_30.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_30.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_30.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_31.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_31.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_31.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_31.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_32.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_32.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_32.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_32.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_33.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_33.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_33.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_33.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_34.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_34.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_34.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_34.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_35.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_35.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_35.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_35.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_36.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_36.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_36.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_36.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_37.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_37.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_37.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_37.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_38.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_38.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_38.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_38.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_39.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_39.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_39.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_39.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_4.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_4.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_4.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_4.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_40.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_40.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_40.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_40.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_41.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_41.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_41.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_41.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_42.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_42.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_42.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_42.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_43.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_43.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_43.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_43.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_44.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_44.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_44.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_44.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_45.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_45.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_45.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_45.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_46.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_46.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_46.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_46.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_47.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_47.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_47.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_47.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_48.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_48.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_48.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_48.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_49.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_49.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_49.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_49.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_5.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_5.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_5.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_5.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_50.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_50.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_50.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_50.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_51.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_51.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_51.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_51.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_6.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_6.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_6.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_6.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_7.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_7.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_7.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_7.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_8.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_8.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_8.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_8.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_9.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_9.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_9.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_9.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_10.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_10.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_10.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_10.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_11.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_11.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_11.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_11.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_12.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_12.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_12.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_12.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_13.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_13.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_13.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_13.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_14.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_14.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_14.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_14.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_15.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_15.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_15.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_15.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_16.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_16.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_16.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_16.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_17.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_17.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_17.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_17.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_18.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_18.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_18.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_18.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_19.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_19.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_19.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_19.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_20.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_20.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_20.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_20.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_21.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_21.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_21.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_21.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_22.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_22.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_22.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_22.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_23.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_23.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_23.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_23.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_24.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_24.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_24.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_24.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_25.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_25.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_25.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_25.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_26.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_26.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_26.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_26.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_27.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_27.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_27.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_27.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_28.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_28.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_28.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_28.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_29.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_29.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_29.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_29.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_30.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_30.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_30.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_30.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_31.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_31.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_31.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_31.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_32.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_32.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_32.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_32.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_33.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_33.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_33.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_33.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_34.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_34.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_34.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_34.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_35.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_35.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_35.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_35.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_36.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_36.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_36.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_36.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_37.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_37.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_37.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_37.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_38.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_38.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_38.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_38.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_39.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_39.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_39.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_39.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_4.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_4.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_4.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_4.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_40.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_40.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_40.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_40.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_41.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_41.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_41.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_41.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_42.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_42.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_42.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_42.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_43.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_43.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_43.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_43.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_44.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_44.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_44.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_44.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_45.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_45.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_45.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_45.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_46.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_46.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_46.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_46.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_47.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_47.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_47.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_47.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_48.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_48.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_48.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_48.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_49.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_49.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_49.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_49.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_5.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_5.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_5.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_5.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_50.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_50.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_50.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_50.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_51.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_51.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_51.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_51.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_6.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_6.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_6.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_6.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_7.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_7.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_7.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_7.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_8.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_8.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_8.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_8.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_9.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_9.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_9.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_9.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_10.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_10.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_10.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_10.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_11.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_11.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_11.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_11.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_12.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_12.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_12.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_12.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_13.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_13.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_13.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_13.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_14.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_14.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_14.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_14.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_15.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_15.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_15.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_15.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_16.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_16.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_16.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_16.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_17.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_17.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_17.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_17.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_18.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_18.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_18.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_18.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_19.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_19.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_19.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_19.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_20.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_20.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_20.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_20.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_21.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_21.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_21.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_21.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_22.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_22.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_22.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_22.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_23.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_23.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_23.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_23.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_24.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_24.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_24.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_24.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_25.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_25.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_25.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_25.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_26.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_26.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_26.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_26.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_27.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_27.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_27.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_27.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_28.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_28.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_28.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_28.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_29.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_29.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_29.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_29.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_30.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_30.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_30.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_30.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_31.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_31.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_31.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_31.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_32.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_32.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_32.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_32.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_33.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_33.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_33.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_33.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_34.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_34.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_34.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_34.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_35.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_35.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_35.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_35.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_36.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_36.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_36.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_36.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_37.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_37.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_37.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_37.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_38.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_38.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_38.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_38.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_39.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_39.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_39.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_39.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_4.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_4.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_4.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_4.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_40.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_40.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_40.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_40.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_41.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_41.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_41.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_41.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_42.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_42.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_42.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_42.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_43.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_43.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_43.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_43.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_44.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_44.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_44.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_44.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_45.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_45.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_45.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_45.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_46.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_46.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_46.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_46.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_47.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_47.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_47.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_47.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_48.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_48.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_48.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_48.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_49.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_49.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_49.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_49.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_5.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_5.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_5.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_5.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_50.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_50.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_50.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_50.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_51.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_51.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_51.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_51.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_6.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_6.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_6.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_6.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_7.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_7.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_7.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_7.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_8.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_8.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_8.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_8.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_9.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_9.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_9.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_9.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_accum_thresh.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_accum_thresh.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_accum_thresh.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_accum_thresh.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_lock.q == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_lock.q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_lock.qe    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_lock.qe &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase0_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase0_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase0_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase0_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase1_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase1_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase1_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase1_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase2_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase2_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase2_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase2_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase3_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase3_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase3_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase3_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_timeout_cyc.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_timeout_cyc.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_timeout_cyc.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_timeout_cyc.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_accum_thresh.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_accum_thresh.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_accum_thresh.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_accum_thresh.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_lock.q == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_lock.q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_lock.qe    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_lock.qe &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase0_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase0_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase0_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase0_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase1_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase1_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase1_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase1_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase2_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase2_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase2_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase2_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase3_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase3_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase3_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase3_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_timeout_cyc.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_timeout_cyc.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_timeout_cyc.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_timeout_cyc.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_accum_thresh.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_accum_thresh.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_accum_thresh.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_accum_thresh.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_lock.q == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_lock.q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_lock.qe    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_lock.qe &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase0_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase0_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase0_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase0_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase1_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase1_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase1_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase1_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase2_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase2_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase2_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase2_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase3_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase3_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase3_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase3_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_timeout_cyc.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_timeout_cyc.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_timeout_cyc.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_timeout_cyc.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_accum_thresh.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_accum_thresh.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_accum_thresh.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_accum_thresh.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_lock.q == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_lock.q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_lock.qe    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_lock.qe &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase0_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase0_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase0_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase0_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase1_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase1_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase1_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase1_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase2_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase2_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase2_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase2_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase3_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase3_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase3_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase3_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_timeout_cyc.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_timeout_cyc.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_timeout_cyc.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_timeout_cyc.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classa.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classa.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classa.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classa.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classb.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classb.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classb.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classb.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classc.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classc.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classc.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classc.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classd.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classd.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classd.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classd.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classa.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classa.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classa.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classa.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classb.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classb.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classb.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classb.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classd.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classd.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classd.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classd.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_4.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_4.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_4.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_4.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_4.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_4.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_4.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_4.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_4.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_4.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_4.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_4.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_4.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_4.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_4.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_4.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timeout_cyc.q == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timeout_cyc.q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timeout_cyc.qe    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timeout_cyc.qe &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_en.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_en.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_en.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_en.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.aon_rst_req_q == top_level_upec.top_earlgrey_2.u_aon_timer_aon.aon_rst_req_q  &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.aon_wkup_req_q    == top_level_upec.top_earlgrey_2.u_aon_timer_aon.aon_wkup_req_q &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.prescale_count_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.prescale_count_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wdog_bark_thold_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wdog_bark_thold_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wdog_bite_thold_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wdog_bite_thold_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wdog_count_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wdog_count_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wdog_enable_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wdog_enable_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wdog_pause_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wdog_pause_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wkup_count_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wkup_count_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wkup_enable_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wkup_enable_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wkup_prescaler_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wkup_prescaler_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wkup_thold_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wkup_thold_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_intr_hw.intr_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_intr_hw.intr_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_intr_state_wdog_timer_expired.q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_intr_state_wdog_timer_expired.q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_intr_state_wdog_timer_expired.qe  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_intr_state_wdog_timer_expired.qe   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_intr_state_wkup_timer_expired.q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_intr_state_wkup_timer_expired.q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_intr_state_wkup_timer_expired.qe  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_intr_state_wkup_timer_expired.qe   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_wdog_regwen.q == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_wdog_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_wdog_regwen.qe    == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_wdog_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_sleep_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_sleep_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_sleep_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_sleep_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_wdog_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_wdog_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_wdog_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_wdog_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_wkup_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_wkup_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_wkup_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_wkup_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_gray_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_sync_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_sync_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_wptr_gray_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_wptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_wptr_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_wptr_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.storage   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.storage    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_gray_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_sync_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_sync_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_wptr_gray_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_wptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_wptr_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_wptr_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.storage   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.storage    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.clk_status   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.clk_status    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.dis_status_q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.dis_status_q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.en_status_q  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.en_status_q   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div2_peri_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div2_peri_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div2_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div2_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div2_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div2_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div4_peri_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div4_peri_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div4_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div4_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div4_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div4_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_peri_cg.gen_generic.u_impl_generic.en_latch == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_peri_cg.gen_generic.u_impl_generic.en_latch  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_aes_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_aes_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_aes_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_aes_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_aes_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_aes_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_hmac_cg.gen_generic.u_impl_generic.en_latch   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_hmac_cg.gen_generic.u_impl_generic.en_latch    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_hmac_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_hmac_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_hmac_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_hmac_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_kmac_cg.gen_generic.u_impl_generic.en_latch   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_kmac_cg.gen_generic.u_impl_generic.en_latch    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_kmac_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_kmac_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_kmac_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_kmac_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_otbn_cg.gen_generic.u_impl_generic.en_latch   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_otbn_cg.gen_generic.u_impl_generic.en_latch    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_otbn_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_otbn_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_otbn_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_otbn_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_usb_peri_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_usb_peri_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_usb_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_usb_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_usb_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_usb_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clkmgr_byp.u_clk_byp_req.u_prim_flop.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clkmgr_byp.u_clk_byp_req.u_prim_flop.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clkmgr_byp.u_rcv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clkmgr_byp.u_rcv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clkmgr_byp.u_rcv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clkmgr_byp.u_rcv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clkmgr_byp.u_send.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clkmgr_byp.u_send.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_cg.i_cg.gen_generic.u_impl_generic.en_latch == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_cg.i_cg.gen_generic.u_impl_generic.en_latch  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div2_cg.i_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div2_cg.i_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div2_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div2_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div2_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div2_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div4_cg.i_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div4_cg.i_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div4_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div4_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div4_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div4_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_main_cg.i_cg.gen_generic.u_impl_generic.en_latch   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_main_cg.i_cg.gen_generic.u_impl_generic.en_latch    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_main_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_main_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_main_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_main_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_no_scan_io_div2_div.gen_div2.step_down_nq  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_no_scan_io_div2_div.gen_div2.step_down_nq   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_no_scan_io_div2_div.gen_div2.u_div2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_no_scan_io_div2_div.gen_div2.u_div2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_no_scan_io_div4_div.clk_int    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_no_scan_io_div4_div.clk_int &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_no_scan_io_div4_div.gen_div.cnt    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_no_scan_io_div4_div.gen_div.cnt &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_no_scan_io_div4_div.step_down_ack_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_no_scan_io_div4_div.step_down_ack_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div2_peri_en.q    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div2_peri_en.q &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div2_peri_en.qe   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div2_peri_en.qe    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div4_peri_en.q    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div4_peri_en.q &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div4_peri_en.qe   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div4_peri_en.qe    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_peri_en.q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_peri_en.q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_peri_en.qe    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_peri_en.qe &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_usb_peri_en.q    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_usb_peri_en.q &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_usb_peri_en.qe   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_usb_peri_en.qe    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_aes_hint.q    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_aes_hint.q &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_aes_hint.qe   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_aes_hint.qe    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_hmac_hint.q   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_hmac_hint.q    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_hmac_hint.qe  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_hmac_hint.qe   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_kmac_hint.q   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_kmac_hint.q    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_kmac_hint.qe  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_kmac_hint.qe   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_otbn_hint.q   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_otbn_hint.q    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_otbn_hint.qe  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_otbn_hint.qe   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_aes_val.q  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_aes_val.q   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_aes_val.qe == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_aes_val.qe  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_hmac_val.q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_hmac_val.q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_hmac_val.qe    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_hmac_val.qe &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_kmac_val.q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_kmac_val.q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_kmac_val.qe    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_kmac_val.qe &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_otbn_val.q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_otbn_val.q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_otbn_val.qe    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_otbn_val.qe &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_extclk_sel.q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_extclk_sel.q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_extclk_sel.qe    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_extclk_sel.qe &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_extclk_sel_regwen.q  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_extclk_sel_regwen.q   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_extclk_sel_regwen.qe == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_extclk_sel_regwen.qe  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_jitter_enable.q  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_jitter_enable.q   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_jitter_enable.qe == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_jitter_enable.qe  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_roots_en_status_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_roots_en_status_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_roots_en_status_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_roots_en_status_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_roots_or_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_roots_or_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_roots_or_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_roots_or_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_usb_cg.i_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_usb_cg.i_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_usb_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_usb_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_usb_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_usb_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_gpio.cio_gpio_en_q  == top_level_upec.top_earlgrey_2.u_gpio.cio_gpio_en_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.cio_gpio_q == top_level_upec.top_earlgrey_2.u_gpio.cio_gpio_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.data_in_q  == top_level_upec.top_earlgrey_2.u_gpio.data_in_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[0].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[0].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[0].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[0].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[0].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[0].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[10].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[10].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[10].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[10].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[10].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[10].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[11].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[11].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[11].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[11].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[11].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[11].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[12].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[12].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[12].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[12].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[12].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[12].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[13].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[13].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[13].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[13].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[13].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[13].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[14].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[14].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[14].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[14].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[14].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[14].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[15].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[15].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[15].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[15].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[15].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[15].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[16].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[16].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[16].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[16].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[16].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[16].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[17].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[17].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[17].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[17].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[17].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[17].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[18].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[18].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[18].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[18].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[18].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[18].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[19].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[19].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[19].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[19].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[19].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[19].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[1].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[1].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[1].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[1].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[1].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[1].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[20].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[20].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[20].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[20].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[20].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[20].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[21].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[21].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[21].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[21].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[21].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[21].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[22].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[22].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[22].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[22].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[22].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[22].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[23].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[23].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[23].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[23].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[23].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[23].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[24].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[24].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[24].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[24].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[24].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[24].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[25].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[25].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[25].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[25].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[25].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[25].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[26].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[26].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[26].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[26].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[26].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[26].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[27].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[27].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[27].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[27].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[27].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[27].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[28].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[28].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[28].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[28].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[28].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[28].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[29].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[29].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[29].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[29].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[29].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[29].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[2].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[2].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[2].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[2].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[2].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[2].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[30].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[30].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[30].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[30].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[30].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[30].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[31].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[31].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[31].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[31].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[31].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[31].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[3].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[3].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[3].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[3].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[3].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[3].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[4].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[4].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[4].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[4].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[4].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[4].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[5].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[5].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[5].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[5].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[5].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[5].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[6].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[6].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[6].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[6].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[6].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[6].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[7].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[7].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[7].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[7].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[7].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[7].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[8].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[8].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[8].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[8].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[8].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[8].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[9].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[9].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[9].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[9].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[9].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[9].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.intr_hw.intr_o == top_level_upec.top_earlgrey_2.u_gpio.intr_hw.intr_o  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_ctrl_en_input_filter.q == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_ctrl_en_input_filter.q  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_ctrl_en_input_filter.qe    == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_ctrl_en_input_filter.qe &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_data_in.q  == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_data_in.q   &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_data_in.qe == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_data_in.qe  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_falling.q == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_falling.q  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_falling.qe    == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_falling.qe &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_lvlhigh.q == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_lvlhigh.q  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_lvlhigh.qe    == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_lvlhigh.qe &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_lvllow.q  == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_lvllow.q   &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_lvllow.qe == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_lvllow.qe  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_rising.q  == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_rising.q   &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_rising.qe == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_rising.qe  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_enable.q  == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_enable.q   &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_enable.qe == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_enable.qe  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_state.q   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_state.q    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_state.qe  == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_state.qe   &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.fmt_watermark_q   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.fmt_watermark_q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_ack_stop.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_ack_stop.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_acq_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_acq_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_fmt_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_fmt_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_fmt_watermark.intr_o  == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_fmt_watermark.intr_o   &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_host_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_host_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_nak.intr_o    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_nak.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_rx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_rx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_rx_watermark.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_rx_watermark.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_scl_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_scl_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_sda_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_sda_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_sda_unstable.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_sda_unstable.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_stretch_timeout.intr_o    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_stretch_timeout.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_trans_complete.intr_o == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_trans_complete.intr_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_tx_empty.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_tx_empty.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_tx_nonempty.intr_o    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_tx_nonempty.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_tx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_tx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.rx_watermark_q    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.rx_watermark_q &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.scl_rx_val    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.scl_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.sda_rx_val    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.sda_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.bit_idx == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.bit_idx  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.bit_index   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.bit_index    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.byte_index  == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.byte_index   &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.host_ack    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.host_ack &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.input_byte  == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.input_byte   &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.no_stop == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.no_stop  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.read_byte   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.read_byte    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.scl_high_cnt    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.scl_high_cnt &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.scl_i_q == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.scl_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.sda_i_q == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.sda_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.start_det   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.start_det    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.state_q == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.state_q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.stop_det    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.stop_det &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.stretch == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.stretch  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.stretch_stop_acq_clr    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.stretch_stop_acq_clr &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.stretch_stop_tx_clr == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.stretch_stop_tx_clr  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.tcount_q    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.tcount_q &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_enablehost.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_enablehost.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_enablehost.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_enablehost.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_enabletarget.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_enabletarget.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_enabletarget.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_enabletarget.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_llpbk.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_llpbk.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_llpbk.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_llpbk.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_fbyte.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_fbyte.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_fbyte.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_fbyte.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_nakok.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_nakok.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_nakok.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_nakok.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_rcont.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_rcont.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_rcont.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_rcont.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_read.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_read.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_read.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_read.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_start.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_start.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_start.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_start.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_stop.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_stop.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_stop.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_stop.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_acqrst.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_acqrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_acqrst.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_acqrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_fmtilvl.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_fmtilvl.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_fmtilvl.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_fmtilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_fmtrst.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_fmtrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_fmtrst.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_fmtrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_rxilvl.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_rxilvl.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_rxilvl.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_rxilvl.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_rxrst.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_rxrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_rxrst.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_rxrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_txrst.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_txrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_txrst.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_txrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_host_timeout_ctrl.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_host_timeout_ctrl.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_host_timeout_ctrl.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_host_timeout_ctrl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_ack_stop.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_ack_stop.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_ack_stop.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_ack_stop.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_acq_overflow.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_acq_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_acq_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_acq_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_fmt_overflow.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_fmt_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_fmt_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_fmt_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_fmt_watermark.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_fmt_watermark.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_fmt_watermark.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_fmt_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_host_timeout.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_host_timeout.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_host_timeout.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_host_timeout.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_nak.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_nak.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_nak.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_nak.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_rx_watermark.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_scl_interference.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_scl_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_scl_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_scl_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_sda_interference.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_sda_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_sda_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_sda_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_sda_unstable.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_sda_unstable.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_sda_unstable.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_sda_unstable.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_stretch_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_stretch_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_stretch_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_stretch_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_trans_complete.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_trans_complete.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_trans_complete.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_trans_complete.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_empty.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_nonempty.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_nonempty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_nonempty.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_nonempty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_ack_stop.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_ack_stop.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_ack_stop.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_ack_stop.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_acq_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_acq_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_acq_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_acq_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_fmt_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_fmt_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_fmt_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_fmt_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_fmt_watermark.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_fmt_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_fmt_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_fmt_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_host_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_host_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_host_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_host_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_nak.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_nak.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_nak.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_nak.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_rx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_rx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_rx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_rx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_rx_watermark.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_rx_watermark.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_rx_watermark.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_rx_watermark.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_scl_interference.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_scl_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_scl_interference.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_scl_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_sda_interference.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_sda_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_sda_interference.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_sda_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_sda_unstable.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_sda_unstable.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_sda_unstable.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_sda_unstable.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_stretch_timeout.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_stretch_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_stretch_timeout.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_stretch_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_trans_complete.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_trans_complete.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_trans_complete.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_trans_complete.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_empty.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_empty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_empty.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_empty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_nonempty.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_nonempty.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_nonempty.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_nonempty.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_sclval.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_sclval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_sclval.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_sclval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_sdaval.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_sdaval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_sdaval.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_sdaval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_txovrden.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_txovrden.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_txovrden.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_txovrden.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_en_addr_acq.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_en_addr_acq.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_en_addr_acq.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_en_addr_acq.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_en_addr_tx.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_en_addr_tx.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_en_addr_tx.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_en_addr_tx.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_stop_acq.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_stop_acq.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_stop_acq.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_stop_acq.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_stop_tx.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_stop_tx.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_stop_tx.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_stop_tx.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_address0.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_address0.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_address0.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_address0.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_address1.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_address1.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_address1.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_address1.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_mask0.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_mask0.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_mask0.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_mask0.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_mask1.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_mask1.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_mask1.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_mask1.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timeout_ctrl_en.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timeout_ctrl_en.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timeout_ctrl_en.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timeout_ctrl_en.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timeout_ctrl_val.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timeout_ctrl_val.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timeout_ctrl_val.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timeout_ctrl_val.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing0_thigh.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing0_thigh.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing0_thigh.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing0_thigh.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing0_tlow.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing0_tlow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing0_tlow.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing0_tlow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing1_t_f.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing1_t_f.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing1_t_f.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing1_t_f.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing1_t_r.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing1_t_r.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing1_t_r.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing1_t_r.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing2_thd_sta.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing2_thd_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing2_thd_sta.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing2_thd_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing2_tsu_sta.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing2_tsu_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing2_tsu_sta.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing2_tsu_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing3_thd_dat.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing3_thd_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing3_thd_dat.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing3_thd_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing3_tsu_dat.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing3_tsu_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing3_tsu_dat.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing3_tsu_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing4_t_buf.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing4_t_buf.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing4_t_buf.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing4_t_buf.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing4_tsu_sto.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing4_tsu_sto.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing4_tsu_sto.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing4_tsu_sto.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_txdata.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_txdata.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_txdata.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_txdata.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.fmt_watermark_q   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.fmt_watermark_q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_ack_stop.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_ack_stop.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_acq_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_acq_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_fmt_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_fmt_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_fmt_watermark.intr_o  == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_fmt_watermark.intr_o   &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_host_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_host_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_nak.intr_o    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_nak.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_rx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_rx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_rx_watermark.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_rx_watermark.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_scl_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_scl_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_sda_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_sda_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_sda_unstable.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_sda_unstable.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_stretch_timeout.intr_o    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_stretch_timeout.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_trans_complete.intr_o == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_trans_complete.intr_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_tx_empty.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_tx_empty.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_tx_nonempty.intr_o    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_tx_nonempty.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_tx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_tx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.rx_watermark_q    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.rx_watermark_q &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.scl_rx_val    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.scl_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.sda_rx_val    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.sda_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.bit_idx == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.bit_idx  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.bit_index   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.bit_index    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.byte_index  == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.byte_index   &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.host_ack    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.host_ack &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.input_byte  == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.input_byte   &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.no_stop == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.no_stop  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.read_byte   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.read_byte    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.scl_high_cnt    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.scl_high_cnt &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.scl_i_q == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.scl_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.sda_i_q == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.sda_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.start_det   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.start_det    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.state_q == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.state_q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.stop_det    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.stop_det &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.stretch == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.stretch  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.stretch_stop_acq_clr    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.stretch_stop_acq_clr &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.stretch_stop_tx_clr == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.stretch_stop_tx_clr  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.tcount_q    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.tcount_q &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_enablehost.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_enablehost.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_enablehost.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_enablehost.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_enabletarget.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_enabletarget.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_enabletarget.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_enabletarget.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_llpbk.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_llpbk.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_llpbk.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_llpbk.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_fbyte.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_fbyte.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_fbyte.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_fbyte.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_nakok.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_nakok.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_nakok.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_nakok.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_rcont.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_rcont.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_rcont.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_rcont.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_read.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_read.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_read.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_read.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_start.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_start.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_start.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_start.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_stop.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_stop.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_stop.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_stop.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_acqrst.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_acqrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_acqrst.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_acqrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_fmtilvl.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_fmtilvl.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_fmtilvl.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_fmtilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_fmtrst.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_fmtrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_fmtrst.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_fmtrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_rxilvl.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_rxilvl.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_rxilvl.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_rxilvl.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_rxrst.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_rxrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_rxrst.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_rxrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_txrst.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_txrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_txrst.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_txrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_host_timeout_ctrl.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_host_timeout_ctrl.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_host_timeout_ctrl.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_host_timeout_ctrl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_ack_stop.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_ack_stop.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_ack_stop.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_ack_stop.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_acq_overflow.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_acq_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_acq_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_acq_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_fmt_overflow.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_fmt_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_fmt_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_fmt_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_fmt_watermark.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_fmt_watermark.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_fmt_watermark.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_fmt_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_host_timeout.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_host_timeout.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_host_timeout.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_host_timeout.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_nak.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_nak.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_nak.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_nak.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_rx_watermark.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_scl_interference.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_scl_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_scl_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_scl_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_sda_interference.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_sda_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_sda_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_sda_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_sda_unstable.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_sda_unstable.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_sda_unstable.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_sda_unstable.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_stretch_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_stretch_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_stretch_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_stretch_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_trans_complete.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_trans_complete.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_trans_complete.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_trans_complete.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_empty.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_nonempty.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_nonempty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_nonempty.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_nonempty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_ack_stop.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_ack_stop.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_ack_stop.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_ack_stop.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_acq_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_acq_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_acq_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_acq_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_fmt_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_fmt_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_fmt_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_fmt_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_fmt_watermark.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_fmt_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_fmt_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_fmt_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_host_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_host_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_host_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_host_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_nak.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_nak.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_nak.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_nak.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_rx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_rx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_rx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_rx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_rx_watermark.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_rx_watermark.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_rx_watermark.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_rx_watermark.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_scl_interference.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_scl_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_scl_interference.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_scl_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_sda_interference.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_sda_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_sda_interference.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_sda_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_sda_unstable.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_sda_unstable.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_sda_unstable.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_sda_unstable.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_stretch_timeout.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_stretch_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_stretch_timeout.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_stretch_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_trans_complete.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_trans_complete.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_trans_complete.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_trans_complete.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_empty.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_empty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_empty.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_empty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_nonempty.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_nonempty.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_nonempty.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_nonempty.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_sclval.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_sclval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_sclval.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_sclval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_sdaval.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_sdaval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_sdaval.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_sdaval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_txovrden.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_txovrden.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_txovrden.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_txovrden.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_en_addr_acq.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_en_addr_acq.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_en_addr_acq.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_en_addr_acq.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_en_addr_tx.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_en_addr_tx.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_en_addr_tx.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_en_addr_tx.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_stop_acq.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_stop_acq.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_stop_acq.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_stop_acq.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_stop_tx.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_stop_tx.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_stop_tx.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_stop_tx.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_address0.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_address0.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_address0.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_address0.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_address1.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_address1.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_address1.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_address1.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_mask0.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_mask0.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_mask0.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_mask0.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_mask1.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_mask1.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_mask1.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_mask1.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timeout_ctrl_en.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timeout_ctrl_en.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timeout_ctrl_en.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timeout_ctrl_en.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timeout_ctrl_val.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timeout_ctrl_val.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timeout_ctrl_val.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timeout_ctrl_val.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing0_thigh.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing0_thigh.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing0_thigh.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing0_thigh.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing0_tlow.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing0_tlow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing0_tlow.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing0_tlow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing1_t_f.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing1_t_f.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing1_t_f.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing1_t_f.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing1_t_r.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing1_t_r.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing1_t_r.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing1_t_r.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing2_thd_sta.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing2_thd_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing2_thd_sta.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing2_thd_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing2_tsu_sta.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing2_tsu_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing2_tsu_sta.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing2_tsu_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing3_thd_dat.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing3_thd_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing3_thd_dat.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing3_thd_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing3_tsu_dat.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing3_tsu_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing3_tsu_dat.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing3_tsu_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing4_t_buf.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing4_t_buf.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing4_t_buf.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing4_t_buf.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing4_tsu_sto.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing4_tsu_sto.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing4_tsu_sto.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing4_tsu_sto.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_txdata.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_txdata.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_txdata.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_txdata.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.fmt_watermark_q   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.fmt_watermark_q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_ack_stop.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_ack_stop.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_acq_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_acq_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_fmt_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_fmt_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_fmt_watermark.intr_o  == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_fmt_watermark.intr_o   &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_host_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_host_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_nak.intr_o    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_nak.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_rx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_rx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_rx_watermark.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_rx_watermark.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_scl_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_scl_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_sda_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_sda_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_sda_unstable.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_sda_unstable.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_stretch_timeout.intr_o    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_stretch_timeout.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_trans_complete.intr_o == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_trans_complete.intr_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_tx_empty.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_tx_empty.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_tx_nonempty.intr_o    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_tx_nonempty.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_tx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_tx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.rx_watermark_q    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.rx_watermark_q &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.scl_rx_val    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.scl_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.sda_rx_val    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.sda_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.bit_idx == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.bit_idx  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.bit_index   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.bit_index    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.byte_index  == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.byte_index   &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.host_ack    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.host_ack &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.input_byte  == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.input_byte   &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.no_stop == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.no_stop  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.read_byte   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.read_byte    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.scl_high_cnt    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.scl_high_cnt &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.scl_i_q == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.scl_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.sda_i_q == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.sda_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.start_det   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.start_det    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.state_q == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.state_q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.stop_det    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.stop_det &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.stretch == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.stretch  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.stretch_stop_acq_clr    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.stretch_stop_acq_clr &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.stretch_stop_tx_clr == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.stretch_stop_tx_clr  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.tcount_q    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.tcount_q &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_enablehost.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_enablehost.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_enablehost.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_enablehost.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_enabletarget.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_enabletarget.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_enabletarget.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_enabletarget.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_llpbk.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_llpbk.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_llpbk.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_llpbk.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_fbyte.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_fbyte.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_fbyte.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_fbyte.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_nakok.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_nakok.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_nakok.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_nakok.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_rcont.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_rcont.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_rcont.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_rcont.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_read.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_read.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_read.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_read.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_start.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_start.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_start.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_start.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_stop.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_stop.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_stop.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_stop.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_acqrst.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_acqrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_acqrst.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_acqrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_fmtilvl.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_fmtilvl.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_fmtilvl.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_fmtilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_fmtrst.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_fmtrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_fmtrst.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_fmtrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_rxilvl.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_rxilvl.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_rxilvl.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_rxilvl.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_rxrst.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_rxrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_rxrst.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_rxrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_txrst.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_txrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_txrst.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_txrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_host_timeout_ctrl.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_host_timeout_ctrl.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_host_timeout_ctrl.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_host_timeout_ctrl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_ack_stop.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_ack_stop.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_ack_stop.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_ack_stop.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_acq_overflow.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_acq_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_acq_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_acq_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_fmt_overflow.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_fmt_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_fmt_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_fmt_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_fmt_watermark.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_fmt_watermark.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_fmt_watermark.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_fmt_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_host_timeout.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_host_timeout.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_host_timeout.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_host_timeout.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_nak.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_nak.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_nak.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_nak.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_rx_watermark.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_scl_interference.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_scl_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_scl_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_scl_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_sda_interference.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_sda_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_sda_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_sda_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_sda_unstable.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_sda_unstable.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_sda_unstable.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_sda_unstable.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_stretch_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_stretch_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_stretch_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_stretch_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_trans_complete.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_trans_complete.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_trans_complete.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_trans_complete.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_empty.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_nonempty.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_nonempty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_nonempty.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_nonempty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_ack_stop.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_ack_stop.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_ack_stop.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_ack_stop.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_acq_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_acq_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_acq_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_acq_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_fmt_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_fmt_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_fmt_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_fmt_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_fmt_watermark.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_fmt_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_fmt_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_fmt_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_host_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_host_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_host_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_host_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_nak.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_nak.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_nak.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_nak.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_rx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_rx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_rx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_rx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_rx_watermark.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_rx_watermark.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_rx_watermark.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_rx_watermark.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_scl_interference.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_scl_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_scl_interference.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_scl_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_sda_interference.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_sda_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_sda_interference.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_sda_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_sda_unstable.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_sda_unstable.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_sda_unstable.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_sda_unstable.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_stretch_timeout.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_stretch_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_stretch_timeout.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_stretch_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_trans_complete.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_trans_complete.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_trans_complete.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_trans_complete.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_empty.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_empty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_empty.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_empty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_nonempty.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_nonempty.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_nonempty.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_nonempty.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_sclval.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_sclval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_sclval.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_sclval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_sdaval.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_sdaval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_sdaval.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_sdaval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_txovrden.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_txovrden.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_txovrden.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_txovrden.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_en_addr_acq.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_en_addr_acq.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_en_addr_acq.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_en_addr_acq.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_en_addr_tx.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_en_addr_tx.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_en_addr_tx.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_en_addr_tx.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_stop_acq.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_stop_acq.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_stop_acq.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_stop_acq.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_stop_tx.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_stop_tx.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_stop_tx.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_stop_tx.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_address0.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_address0.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_address0.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_address0.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_address1.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_address1.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_address1.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_address1.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_mask0.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_mask0.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_mask0.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_mask0.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_mask1.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_mask1.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_mask1.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_mask1.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timeout_ctrl_en.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timeout_ctrl_en.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timeout_ctrl_en.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timeout_ctrl_en.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timeout_ctrl_val.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timeout_ctrl_val.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timeout_ctrl_val.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timeout_ctrl_val.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing0_thigh.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing0_thigh.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing0_thigh.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing0_thigh.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing0_tlow.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing0_tlow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing0_tlow.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing0_tlow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing1_t_f.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing1_t_f.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing1_t_f.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing1_t_f.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing1_t_r.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing1_t_r.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing1_t_r.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing1_t_r.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing2_thd_sta.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing2_thd_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing2_thd_sta.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing2_thd_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing2_tsu_sta.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing2_tsu_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing2_tsu_sta.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing2_tsu_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing3_thd_dat.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing3_thd_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing3_thd_dat.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing3_thd_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing3_tsu_dat.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing3_tsu_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing3_tsu_dat.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing3_tsu_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing4_t_buf.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing4_t_buf.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing4_t_buf.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing4_t_buf.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing4_tsu_sto.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing4_tsu_sto.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing4_tsu_sto.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing4_tsu_sto.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_txdata.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_txdata.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_txdata.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_txdata.qe   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.fatal_bus_integ_error_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.fatal_bus_integ_error_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.fatal_prog_error_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.fatal_prog_error_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.fatal_state_error_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.fatal_state_error_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.flash_rma_error_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.flash_rma_error_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_set_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_set_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.ping_set_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.state_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.state_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_set_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_set_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_test_set_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_test_set_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.ping_set_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.ping_set_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.state_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.state_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.level_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.level_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.level_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.level_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_prim_generic_flop.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_prim_generic_flop.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.alert_set_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.alert_set_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.alert_test_set_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.alert_test_set_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.ping_set_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.ping_set_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.state_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.state_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ack.level_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ack.level_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ping.level_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ping.level_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_prim_generic_flop.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_prim_generic_flop.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_done_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_done_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_idle_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_idle_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.otp_part_error_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.otp_part_error_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.otp_test_ctrl_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.otp_test_ctrl_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.sw_claim_transition_if_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.sw_claim_transition_if_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.tap_claim_transition_if_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.tap_claim_transition_if_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.token_invalid_error_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.token_invalid_error_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.trans_cnt_oflw_error_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.trans_cnt_oflw_error_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.trans_invalid_error_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.trans_invalid_error_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.trans_success_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.trans_success_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.transition_target_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.transition_target_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.transition_token_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.transition_token_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.address_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.address_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.data_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.data_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.dr_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.dr_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.error_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.error_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_gray_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_sync_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_sync_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_wptr_gray_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_wptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_wptr_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_wptr_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.storage  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.storage   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.storage == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.storage  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.bypass_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.bypass_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.dtmcs_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.dtmcs_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.idcode_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.idcode_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.jtag_ir_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.jtag_ir_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.jtag_ir_shift_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.jtag_ir_shift_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.tap_state_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.tap_state_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.td_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.td_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.tdo_oe_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.tdo_oe_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.state_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.state_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.lc_state_valid_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.lc_state_valid_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_cnt_regs.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_cnt_regs.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_fsm_state_regs.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_fsm_state_regs.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_id_state_regs.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_id_state_regs.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_flo_keymgr_div.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_flo_keymgr_div.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_cpu_en.u_prim_flop.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_cpu_en.u_prim_flop.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_creator_seed_sw_rw_en.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_creator_seed_sw_rw_en.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_dft_en.u_prim_flop.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_dft_en.u_prim_flop.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_escalate_en.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_escalate_en.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_hw_debug_en.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_hw_debug_en.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_iso_part_sw_rd_en.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_iso_part_sw_rd_en.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_iso_part_sw_wr_en.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_iso_part_sw_wr_en.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_keymgr_en.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_keymgr_en.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_nvm_debug_en.u_prim_flop.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_nvm_debug_en.u_prim_flop.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_owner_seed_sw_rw_en.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_owner_seed_sw_rw_en.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_seed_hw_rd_en.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_seed_hw_rd_en.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_test_or_rma.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_test_or_rma.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_check_byp_en.u_prim_flop.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_check_byp_en.u_prim_flop.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_clk_byp_req.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_clk_byp_req.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_flash_rma_req.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_flash_rma_req.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_clk_byp_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_clk_byp_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_clk_byp_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_clk_byp_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_flash_rma_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_flash_rma_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_flash_rma_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_flash_rma_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_state_regs.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_state_regs.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.hashed_token_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.hashed_token_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.token_hash_ack_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.token_hash_ack_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.token_hash_err_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.token_hash_err_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.gen_data_reg.data_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.gen_data_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.dst_ack_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.dst_ack_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.dst_fsm_cs  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.dst_fsm_cs   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.src_fsm_cs  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.src_fsm_cs   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.src_req_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.src_req_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.dst_ack_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.dst_ack_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.dst_fsm_cs == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.dst_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.src_fsm_cs == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.src_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.src_req_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.src_req_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_state_regs.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_state_regs.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver1.state_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver1.state_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver1.u_decode_esc.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver1.u_decode_esc.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver1.u_decode_esc.level_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver1.u_decode_esc.level_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver1.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver1.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver2.state_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver2.state_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver2.u_decode_esc.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver2.u_decode_esc.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver2.u_decode_esc.level_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver2.u_decode_esc.level_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver2.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver2.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_flop_2sync_init.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_flop_2sync_init.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_flop_2sync_init.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_flop_2sync_init.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.intg_err_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.intg_err_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_tap_tlul_host.g_multiple_reqs.source_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_tap_tlul_host.g_multiple_reqs.source_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_tap_tlul_host.intg_err_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_tap_tlul_host.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_tap_tlul_host.outstanding_reqs_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_tap_tlul_host.outstanding_reqs_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.fatal_check_error_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.fatal_check_error_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.fatal_macro_error_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.fatal_macro_error_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.pending_tlul_error_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.pending_tlul_error_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.tlul_addr_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.tlul_addr_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.pending_tlul_error_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.pending_tlul_error_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.tlul_addr_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.tlul_addr_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.cnt_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.cnt_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.dout_gate_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.dout_gate_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.cnt_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.cnt_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.dout_gate_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.dout_gate_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.cnt_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.cnt_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.dout_gate_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.dout_gate_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.cnt_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.cnt_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.dout_gate_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.dout_gate_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.cnt_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.cnt_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.dout_gate_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.dout_gate_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.error_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.error_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_otp_ctrl_ecc_reg.data_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_otp_ctrl_ecc_reg.data_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.interrupt_triggers_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.interrupt_triggers_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.otp_idle_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.otp_idle_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.pwr_otp_rsp_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.pwr_otp_rsp_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.tlul_oob_err_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.tlul_oob_err_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_edn_arb.gen_normal_case.prio_mask_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_edn_arb.gen_normal_case.prio_mask_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_intr_esc0.intr_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_intr_esc0.intr_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_intr_esc1.intr_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_intr_esc1.intr_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.addr_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.addr_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.cnt_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.err_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.err_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.rdata_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.rdata_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.size_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.size_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_rdata_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_rdata_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_regfile_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_regfile_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_rvalid_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_rvalid_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.addr_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.addr_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rdata_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.req_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.req_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rerror_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rerror_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rvalid_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rvalid_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rvalid_sram_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rvalid_sram_q    &&
        //top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.mem    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.mem &&
        //top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.rdata_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.rdata_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.wdata_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.wdata_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.wmask_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.wmask_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.write_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.write_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_state_regs.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_state_regs.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.intg_error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.intg_error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.valid_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.valid_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.wdata_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.wdata_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_arb.gen_normal_case.prio_mask_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_arb.gen_normal_case.prio_mask_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_dai.base_sel_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_dai.base_sel_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_dai.cnt_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_dai.cnt_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_dai.data_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_dai.data_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_dai.error_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_dai.error_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_dai.u_state_regs.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_dai.u_state_regs.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.edn_req_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.edn_req_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.entropy_cnt_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.entropy_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.key_out_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.key_out_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.nonce_out_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.nonce_out_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.seed_cnt_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.seed_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.seed_valid_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.seed_valid_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.u_req_arb.gen_normal_case.prio_mask_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.u_req_arb.gen_normal_case.prio_mask_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.u_state_regs.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.u_state_regs.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lci.cnt_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lci.cnt_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lci.error_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lci.error_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lci.u_state_regs.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lci.u_state_regs.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.chk_timeout_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.chk_timeout_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.cnsty_chk_req_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.cnsty_chk_req_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.cnsty_chk_trig_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.cnsty_chk_trig_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[0].u_prim_flop_cnsty_cnt.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[0].u_prim_flop_cnsty_cnt.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[0].u_prim_flop_integ_cnt.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[0].u_prim_flop_integ_cnt.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[1].u_prim_flop_cnsty_cnt.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[1].u_prim_flop_cnsty_cnt.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[1].u_prim_flop_integ_cnt.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[1].u_prim_flop_integ_cnt.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.cnt_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.perturbed_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.perturbed_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.lfsr_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.lfsr_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.cnt_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.perturbed_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.perturbed_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.lfsr_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.lfsr_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.integ_chk_req_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.integ_chk_req_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.integ_chk_trig_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.integ_chk_trig_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.reseed_timer_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.reseed_timer_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_init_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_init_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_init_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_init_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.fips_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.fips_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.clr_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.clr_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.data_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.data_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.depth_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.depth_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_check_byp_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_check_byp_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_check_byp_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_check_byp_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_creator_seed_sw_rw_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_creator_seed_sw_rw_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_creator_seed_sw_rw_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_creator_seed_sw_rw_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_dft_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_dft_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_dft_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_dft_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_seed_hw_rd_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_seed_hw_rd_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_seed_hw_rd_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_seed_hw_rd_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_regwen.q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_regwen.qe    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_timeout.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_timeout.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_timeout.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_timeout.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_trigger_regwen.q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_trigger_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_trigger_regwen.qe    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_trigger_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_consistency_check_period.q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_consistency_check_period.q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_consistency_check_period.qe    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_consistency_check_period.qe &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_creator_sw_cfg_read_lock.q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_creator_sw_cfg_read_lock.q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_creator_sw_cfg_read_lock.qe    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_creator_sw_cfg_read_lock.qe &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_address.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_address.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_address.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_address.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_wdata_0.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_wdata_0.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_wdata_0.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_wdata_0.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_wdata_1.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_wdata_1.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_wdata_1.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_wdata_1.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_integrity_check_period.q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_integrity_check_period.q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_integrity_check_period.qe  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_integrity_check_period.qe   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_enable_otp_error.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_enable_otp_error.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_enable_otp_error.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_enable_otp_error.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_enable_otp_operation_done.q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_enable_otp_operation_done.q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_enable_otp_operation_done.qe  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_enable_otp_operation_done.qe   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_state_otp_error.q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_state_otp_error.q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_state_otp_error.qe    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_state_otp_error.qe &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_state_otp_operation_done.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_state_otp_operation_done.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_state_otp_operation_done.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_state_otp_operation_done.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_owner_sw_cfg_read_lock.q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_owner_sw_cfg_read_lock.q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_owner_sw_cfg_read_lock.qe  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_owner_sw_cfg_read_lock.qe   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.dev_select_outstanding  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.dev_select_outstanding   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.err_resp.err_opcode == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.err_resp.err_opcode  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.err_resp.err_req_pending    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.err_resp.err_req_pending &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.err_resp.err_rsp_pending    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.err_resp.err_rsp_pending &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.err_resp.err_size   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.err_resp.err_size    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.err_resp.err_source == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.err_resp.err_source  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.num_req_outstanding == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.num_req_outstanding  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.cnt_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.data_shadow_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.data_shadow_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.data_state_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.data_state_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.digest_mode_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.digest_mode_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.digest_state_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.digest_state_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.idx_state_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.idx_state_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.key_state_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.key_state_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.u_state_regs.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.u_state_regs.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.valid_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.valid_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl_mtx.gen_normal_case.prio_mask_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl_mtx.gen_normal_case.prio_mask_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.intg_error_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.intg_error_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.alert_set_q == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.alert_set_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.ping_set_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.state_q == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.state_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.bit_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.bit_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.clk_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.clk_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.complete_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.complete_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.complete_q2    == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.complete_q2 &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.data_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.data_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.len_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.len_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.pcl_int_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.pcl_int_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.polarity_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.polarity_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.prediv_q   == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.prediv_q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.rep_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.rep_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.reps_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.reps_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.bit_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.bit_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.clk_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.clk_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.complete_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.complete_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.complete_q2    == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.complete_q2 &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.data_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.data_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.len_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.len_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.pcl_int_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.pcl_int_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.polarity_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.polarity_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.prediv_q   == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.prediv_q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.rep_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.rep_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.reps_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.reps_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.intr_hw_done_ch0.intr_o  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.intr_hw_done_ch0.intr_o   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.intr_hw_done_ch1.intr_o  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.intr_hw_done_ch1.intr_o   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.intg_err_q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_enable_ch0.q   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_enable_ch0.q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_enable_ch0.qe  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_enable_ch0.qe   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_enable_ch1.q   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_enable_ch1.q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_enable_ch1.qe  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_enable_ch1.qe   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_polarity_ch0.q == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_polarity_ch0.q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_polarity_ch0.qe    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_polarity_ch0.qe &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_polarity_ch1.q == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_polarity_ch1.q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_polarity_ch1.qe    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_polarity_ch1.qe &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch0_0.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch0_0.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch0_0.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch0_0.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch0_1.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch0_1.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch0_1.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch0_1.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch1_0.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch1_0.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch1_0.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch1_0.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch1_1.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch1_1.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch1_1.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch1_1.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_enable_done_ch0.q  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_enable_done_ch0.q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_enable_done_ch0.qe == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_enable_done_ch0.qe  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_enable_done_ch1.q  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_enable_done_ch1.q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_enable_done_ch1.qe == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_enable_done_ch1.qe  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_state_done_ch0.q   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_state_done_ch0.q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_state_done_ch0.qe  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_state_done_ch0.qe   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_state_done_ch1.q   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_state_done_ch1.q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_state_done_ch1.qe  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_state_done_ch1.qe   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_prediv_ch0.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_prediv_ch0.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_prediv_ch0.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_prediv_ch0.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_prediv_ch1.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_prediv_ch1.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_prediv_ch1.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_prediv_ch1.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_len_ch0.q  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_len_ch0.q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_len_ch0.qe == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_len_ch0.qe  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_len_ch1.q  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_len_ch1.q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_len_ch1.qe == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_len_ch1.qe  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_reps_ch0.q == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_reps_ch0.q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_reps_ch0.qe    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_reps_ch0.qe &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_reps_ch1.q == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_reps_ch1.q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_reps_ch1.qe    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_reps_ch1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_oe_retreg_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_oe_retreg_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_out_retreg_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_out_retreg_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_pad_attr_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_pad_attr_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.alert_set_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.ping_set_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.state_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.state_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_oe_retreg_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_oe_retreg_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_out_retreg_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_out_retreg_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_pad_attr_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_pad_attr_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.sleep_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.sleep_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.dft_strap_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.dft_strap_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.dft_strap_valid_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.dft_strap_valid_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.tap_strap_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.tap_strap_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_dft.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_dft.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_dft.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_dft.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_rv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_rv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_rv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_rv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_0.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_0.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_0.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_1.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_1.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_1.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_10.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_10.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_10.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_10.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_11.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_11.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_11.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_11.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_12.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_12.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_12.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_12.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_13.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_13.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_13.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_13.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_14.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_14.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_14.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_14.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_15.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_15.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_15.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_15.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_16.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_16.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_16.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_16.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_17.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_17.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_17.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_17.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_18.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_18.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_18.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_18.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_19.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_19.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_19.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_19.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_2.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_2.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_2.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_20.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_20.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_20.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_20.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_21.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_21.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_21.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_21.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_22.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_22.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_22.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_22.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_23.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_23.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_23.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_23.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_3.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_3.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_3.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_4.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_4.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_4.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_5.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_5.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_5.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_6.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_6.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_6.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_6.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_7.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_7.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_7.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_7.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_8.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_8.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_8.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_8.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_9.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_9.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_9.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_9.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_10.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_10.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_10.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_10.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_11.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_11.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_11.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_11.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_12.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_12.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_12.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_12.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_13.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_13.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_13.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_13.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_14.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_14.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_14.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_14.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_15.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_15.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_15.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_15.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_16.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_16.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_16.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_16.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_17.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_17.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_17.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_17.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_18.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_18.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_18.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_18.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_19.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_19.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_19.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_19.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_20.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_20.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_20.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_20.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_21.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_21.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_21.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_21.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_22.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_22.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_22.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_22.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_23.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_23.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_23.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_23.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_8.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_8.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_8.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_8.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_9.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_9.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_9.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_9.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_0.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_0.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_0.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_1.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_1.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_1.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_10.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_10.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_10.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_10.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_11.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_11.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_11.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_11.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_12.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_12.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_12.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_12.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_13.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_13.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_13.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_13.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_14.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_14.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_14.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_14.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_15.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_15.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_15.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_15.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_16.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_16.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_16.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_16.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_17.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_17.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_17.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_17.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_18.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_18.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_18.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_18.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_19.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_19.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_19.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_19.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_2.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_2.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_2.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_20.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_20.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_20.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_20.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_21.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_21.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_21.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_21.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_22.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_22.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_22.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_22.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_23.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_23.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_23.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_23.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_3.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_3.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_3.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_4.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_4.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_4.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_5.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_5.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_5.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_6.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_6.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_6.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_6.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_7.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_7.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_7.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_7.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_8.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_8.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_8.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_8.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_9.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_9.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_9.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_9.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_10.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_10.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_10.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_10.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_11.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_11.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_11.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_11.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_12.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_12.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_12.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_12.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_13.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_13.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_13.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_13.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_14.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_14.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_14.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_14.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_15.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_15.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_15.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_15.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_16.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_16.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_16.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_16.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_17.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_17.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_17.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_17.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_18.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_18.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_18.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_18.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_19.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_19.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_19.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_19.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_20.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_20.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_20.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_20.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_21.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_21.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_21.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_21.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_22.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_22.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_22.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_22.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_23.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_23.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_23.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_23.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_8.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_8.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_8.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_8.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_9.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_9.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_9.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_9.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_0.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_0.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_0.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_1.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_1.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_1.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_10.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_10.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_10.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_10.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_11.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_11.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_11.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_11.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_12.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_12.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_12.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_12.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_13.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_13.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_13.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_13.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_14.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_14.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_14.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_14.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_15.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_15.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_15.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_15.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_16.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_16.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_16.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_16.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_17.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_17.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_17.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_17.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_18.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_18.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_18.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_18.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_19.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_19.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_19.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_19.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_2.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_2.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_2.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_20.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_20.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_20.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_20.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_21.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_21.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_21.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_21.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_22.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_22.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_22.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_22.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_23.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_23.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_23.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_23.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_3.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_3.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_3.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_4.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_4.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_4.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_5.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_5.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_5.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_6.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_6.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_6.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_6.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_7.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_7.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_7.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_7.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_8.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_8.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_8.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_8.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_9.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_9.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_9.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_9.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_0.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_0.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_0.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_1.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_1.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_1.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_10.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_10.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_10.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_10.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_11.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_11.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_11.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_11.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_12.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_12.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_12.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_12.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_13.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_13.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_13.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_13.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_14.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_14.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_14.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_14.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_15.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_15.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_15.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_15.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_16.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_16.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_16.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_16.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_17.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_17.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_17.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_17.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_18.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_18.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_18.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_18.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_19.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_19.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_19.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_19.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_2.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_2.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_2.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_20.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_20.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_20.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_20.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_21.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_21.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_21.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_21.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_22.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_22.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_22.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_22.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_23.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_23.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_23.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_23.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_24.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_24.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_24.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_24.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_25.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_25.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_25.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_25.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_26.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_26.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_26.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_26.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_27.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_27.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_27.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_27.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_28.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_28.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_28.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_28.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_29.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_29.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_29.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_29.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_3.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_3.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_3.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_30.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_30.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_30.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_30.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_31.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_31.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_31.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_31.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_32.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_32.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_32.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_32.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_33.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_33.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_33.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_33.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_34.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_34.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_34.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_34.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_35.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_35.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_35.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_35.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_36.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_36.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_36.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_36.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_37.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_37.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_37.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_37.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_38.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_38.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_38.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_38.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_39.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_39.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_39.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_39.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_4.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_4.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_4.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_40.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_40.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_40.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_40.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_41.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_41.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_41.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_41.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_42.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_42.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_42.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_42.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_43.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_43.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_43.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_43.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_44.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_44.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_44.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_44.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_45.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_45.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_45.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_45.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_46.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_46.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_46.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_46.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_5.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_5.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_5.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_6.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_6.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_6.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_6.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_7.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_7.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_7.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_7.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_8.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_8.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_8.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_8.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_9.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_9.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_9.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_9.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_0.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_0.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_0.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_0.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_1.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_1.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_1.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_1.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_10.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_10.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_10.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_10.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_11.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_11.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_11.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_11.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_12.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_12.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_12.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_12.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_13.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_13.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_13.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_13.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_14.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_14.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_14.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_14.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_15.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_15.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_15.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_15.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_16.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_16.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_16.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_16.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_17.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_17.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_17.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_17.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_18.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_18.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_18.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_18.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_19.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_19.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_19.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_19.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_2.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_2.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_2.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_2.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_20.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_20.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_20.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_20.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_21.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_21.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_21.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_21.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_22.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_22.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_22.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_22.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_23.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_23.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_23.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_23.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_24.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_24.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_24.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_24.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_25.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_25.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_25.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_25.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_26.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_26.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_26.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_26.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_27.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_27.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_27.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_27.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_28.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_28.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_28.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_28.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_29.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_29.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_29.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_29.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_3.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_3.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_3.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_3.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_30.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_30.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_30.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_30.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_31.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_31.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_31.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_31.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_32.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_32.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_32.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_32.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_33.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_33.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_33.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_33.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_34.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_34.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_34.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_34.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_35.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_35.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_35.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_35.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_36.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_36.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_36.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_36.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_37.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_37.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_37.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_37.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_38.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_38.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_38.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_38.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_39.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_39.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_39.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_39.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_4.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_4.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_4.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_4.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_40.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_40.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_40.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_40.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_41.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_41.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_41.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_41.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_42.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_42.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_42.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_42.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_43.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_43.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_43.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_43.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_44.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_44.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_44.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_44.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_45.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_45.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_45.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_45.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_46.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_46.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_46.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_46.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_5.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_5.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_5.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_5.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_6.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_6.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_6.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_6.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_7.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_7.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_7.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_7.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_8.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_8.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_8.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_8.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_9.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_9.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_9.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_9.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_0.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_0.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_0.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_1.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_1.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_1.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_10.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_10.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_10.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_10.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_11.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_11.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_11.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_11.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_12.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_12.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_12.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_12.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_13.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_13.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_13.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_13.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_14.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_14.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_14.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_14.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_15.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_15.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_15.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_15.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_16.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_16.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_16.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_16.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_17.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_17.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_17.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_17.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_18.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_18.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_18.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_18.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_19.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_19.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_19.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_19.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_2.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_2.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_2.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_20.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_20.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_20.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_20.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_21.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_21.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_21.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_21.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_22.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_22.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_22.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_22.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_23.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_23.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_23.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_23.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_24.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_24.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_24.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_24.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_25.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_25.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_25.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_25.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_26.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_26.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_26.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_26.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_27.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_27.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_27.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_27.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_28.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_28.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_28.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_28.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_29.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_29.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_29.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_29.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_3.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_3.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_3.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_30.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_30.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_30.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_30.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_31.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_31.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_31.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_31.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_32.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_32.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_32.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_32.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_33.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_33.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_33.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_33.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_34.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_34.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_34.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_34.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_35.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_35.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_35.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_35.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_36.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_36.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_36.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_36.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_37.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_37.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_37.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_37.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_38.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_38.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_38.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_38.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_39.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_39.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_39.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_39.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_4.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_4.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_4.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_40.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_40.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_40.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_40.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_41.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_41.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_41.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_41.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_42.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_42.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_42.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_42.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_43.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_43.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_43.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_43.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_44.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_44.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_44.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_44.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_45.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_45.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_45.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_45.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_46.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_46.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_46.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_46.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_5.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_5.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_5.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_6.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_6.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_6.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_6.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_7.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_7.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_7.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_7.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_8.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_8.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_8.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_8.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_9.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_9.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_9.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_9.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_10.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_10.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_10.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_10.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_11.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_11.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_11.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_11.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_12.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_12.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_12.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_12.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_13.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_13.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_13.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_13.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_14.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_14.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_14.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_14.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_15.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_15.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_15.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_15.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_16.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_16.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_16.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_16.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_17.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_17.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_17.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_17.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_18.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_18.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_18.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_18.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_19.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_19.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_19.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_19.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_20.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_20.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_20.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_20.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_21.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_21.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_21.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_21.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_22.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_22.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_22.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_22.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_23.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_23.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_23.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_23.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_24.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_24.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_24.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_24.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_25.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_25.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_25.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_25.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_26.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_26.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_26.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_26.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_27.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_27.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_27.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_27.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_28.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_28.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_28.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_28.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_29.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_29.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_29.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_29.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_30.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_30.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_30.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_30.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_31.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_31.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_31.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_31.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_32.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_32.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_32.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_32.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_33.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_33.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_33.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_33.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_34.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_34.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_34.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_34.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_35.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_35.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_35.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_35.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_36.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_36.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_36.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_36.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_37.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_37.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_37.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_37.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_38.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_38.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_38.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_38.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_39.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_39.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_39.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_39.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_40.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_40.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_40.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_40.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_41.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_41.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_41.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_41.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_42.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_42.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_42.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_42.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_43.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_43.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_43.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_43.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_44.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_44.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_44.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_44.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_45.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_45.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_45.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_45.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_46.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_46.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_46.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_46.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_8.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_8.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_8.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_8.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_9.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_9.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_9.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_9.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_0.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_0.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_0.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_1.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_1.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_1.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_10.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_10.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_10.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_10.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_11.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_11.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_11.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_11.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_12.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_12.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_12.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_12.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_13.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_13.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_13.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_13.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_14.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_14.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_14.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_14.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_15.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_15.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_15.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_15.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_16.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_16.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_16.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_16.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_17.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_17.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_17.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_17.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_18.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_18.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_18.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_18.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_19.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_19.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_19.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_19.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_2.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_2.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_2.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_20.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_20.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_20.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_20.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_21.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_21.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_21.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_21.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_22.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_22.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_22.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_22.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_23.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_23.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_23.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_23.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_24.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_24.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_24.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_24.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_25.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_25.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_25.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_25.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_26.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_26.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_26.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_26.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_27.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_27.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_27.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_27.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_28.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_28.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_28.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_28.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_29.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_29.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_29.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_29.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_3.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_3.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_3.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_30.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_30.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_30.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_30.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_31.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_31.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_31.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_31.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_32.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_32.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_32.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_32.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_33.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_33.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_33.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_33.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_34.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_34.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_34.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_34.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_35.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_35.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_35.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_35.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_36.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_36.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_36.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_36.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_37.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_37.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_37.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_37.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_38.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_38.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_38.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_38.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_39.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_39.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_39.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_39.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_4.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_4.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_4.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_40.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_40.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_40.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_40.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_41.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_41.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_41.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_41.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_42.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_42.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_42.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_42.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_43.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_43.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_43.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_43.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_44.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_44.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_44.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_44.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_45.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_45.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_45.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_45.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_46.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_46.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_46.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_46.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_5.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_5.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_5.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_6.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_6.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_6.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_6.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_7.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_7.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_7.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_7.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_8.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_8.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_8.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_8.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_9.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_9.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_9.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_9.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_10.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_10.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_10.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_10.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_11.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_11.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_11.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_11.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_12.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_12.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_12.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_12.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_13.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_13.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_13.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_13.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_14.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_14.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_14.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_14.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_15.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_15.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_15.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_15.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_16.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_16.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_16.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_16.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_17.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_17.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_17.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_17.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_18.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_18.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_18.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_18.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_19.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_19.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_19.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_19.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_20.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_20.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_20.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_20.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_21.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_21.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_21.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_21.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_22.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_22.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_22.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_22.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_23.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_23.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_23.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_23.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_24.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_24.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_24.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_24.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_25.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_25.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_25.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_25.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_26.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_26.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_26.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_26.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_27.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_27.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_27.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_27.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_28.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_28.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_28.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_28.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_29.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_29.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_29.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_29.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_30.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_30.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_30.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_30.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_31.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_31.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_31.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_31.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_32.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_32.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_32.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_32.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_33.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_33.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_33.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_33.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_34.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_34.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_34.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_34.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_35.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_35.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_35.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_35.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_36.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_36.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_36.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_36.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_37.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_37.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_37.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_37.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_38.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_38.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_38.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_38.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_39.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_39.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_39.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_39.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_40.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_40.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_40.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_40.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_41.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_41.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_41.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_41.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_42.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_42.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_42.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_42.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_43.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_43.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_43.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_43.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_44.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_44.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_44.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_44.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_45.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_45.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_45.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_45.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_46.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_46.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_46.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_46.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_8.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_8.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_8.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_8.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_9.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_9.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_9.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_9.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_0.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_0.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_0.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_0.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_1.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_1.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_1.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_1.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_10.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_10.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_10.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_10.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_11.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_11.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_11.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_11.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_12.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_12.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_12.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_12.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_13.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_13.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_13.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_13.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_14.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_14.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_14.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_14.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_15.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_15.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_15.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_15.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_16.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_16.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_16.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_16.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_17.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_17.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_17.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_17.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_18.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_18.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_18.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_18.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_19.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_19.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_19.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_19.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_2.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_2.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_2.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_2.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_20.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_20.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_20.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_20.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_21.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_21.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_21.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_21.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_22.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_22.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_22.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_22.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_23.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_23.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_23.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_23.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_24.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_24.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_24.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_24.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_25.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_25.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_25.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_25.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_26.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_26.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_26.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_26.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_27.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_27.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_27.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_27.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_28.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_28.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_28.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_28.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_29.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_29.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_29.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_29.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_3.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_3.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_3.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_3.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_30.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_30.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_30.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_30.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_31.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_31.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_31.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_31.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_4.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_4.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_4.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_4.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_5.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_5.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_5.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_5.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_6.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_6.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_6.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_6.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_7.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_7.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_7.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_7.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_8.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_8.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_8.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_8.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_9.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_9.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_9.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_9.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_32.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_32.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_32.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_32.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_33.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_33.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_33.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_33.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_34.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_34.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_34.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_34.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_35.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_35.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_35.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_35.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_36.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_36.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_36.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_36.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_37.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_37.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_37.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_37.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_38.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_38.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_38.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_38.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_39.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_39.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_39.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_39.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_40.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_40.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_40.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_40.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_41.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_41.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_41.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_41.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_42.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_42.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_42.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_42.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_43.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_43.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_43.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_43.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_44.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_44.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_44.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_44.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_45.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_45.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_45.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_45.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_46.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_46.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_46.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_46.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_10.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_10.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_10.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_10.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_11.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_11.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_11.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_11.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_12.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_12.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_12.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_12.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_13.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_13.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_13.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_13.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_14.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_14.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_14.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_14.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_15.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_15.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_15.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_15.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_16.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_16.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_16.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_16.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_17.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_17.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_17.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_17.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_18.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_18.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_18.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_18.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_19.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_19.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_19.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_19.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_20.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_20.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_20.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_20.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_21.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_21.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_21.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_21.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_22.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_22.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_22.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_22.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_23.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_23.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_23.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_23.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_24.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_24.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_24.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_24.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_25.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_25.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_25.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_25.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_26.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_26.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_26.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_26.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_27.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_27.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_27.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_27.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_28.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_28.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_28.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_28.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_29.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_29.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_29.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_29.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_30.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_30.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_30.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_30.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_31.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_31.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_31.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_31.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_32.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_32.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_32.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_32.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_33.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_33.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_33.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_33.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_34.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_34.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_34.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_34.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_35.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_35.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_35.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_35.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_36.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_36.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_36.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_36.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_37.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_37.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_37.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_37.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_38.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_38.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_38.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_38.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_39.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_39.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_39.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_39.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_40.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_40.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_40.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_40.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_41.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_41.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_41.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_41.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_42.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_42.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_42.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_42.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_43.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_43.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_43.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_43.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_44.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_44.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_44.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_44.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_45.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_45.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_45.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_45.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_46.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_46.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_46.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_46.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_47.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_47.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_47.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_47.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_48.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_48.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_48.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_48.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_49.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_49.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_49.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_49.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_50.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_50.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_50.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_50.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_51.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_51.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_51.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_51.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_52.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_52.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_52.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_52.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_53.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_53.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_53.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_53.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_54.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_54.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_54.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_54.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_8.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_8.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_8.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_8.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_9.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_9.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_9.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_9.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_0.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_0.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_0.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_1.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_1.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_1.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_10.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_10.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_10.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_10.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_11.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_11.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_11.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_11.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_12.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_12.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_12.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_12.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_13.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_13.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_13.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_13.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_14.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_14.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_14.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_14.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_15.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_15.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_15.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_15.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_16.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_16.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_16.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_16.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_17.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_17.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_17.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_17.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_18.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_18.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_18.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_18.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_19.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_19.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_19.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_19.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_2.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_2.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_2.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_20.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_20.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_20.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_20.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_21.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_21.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_21.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_21.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_22.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_22.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_22.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_22.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_23.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_23.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_23.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_23.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_24.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_24.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_24.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_24.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_25.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_25.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_25.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_25.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_26.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_26.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_26.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_26.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_27.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_27.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_27.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_27.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_28.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_28.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_28.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_28.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_29.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_29.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_29.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_29.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_3.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_3.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_3.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_30.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_30.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_30.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_30.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_31.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_31.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_31.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_31.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_32.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_32.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_32.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_32.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_33.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_33.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_33.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_33.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_34.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_34.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_34.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_34.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_35.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_35.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_35.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_35.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_36.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_36.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_36.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_36.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_37.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_37.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_37.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_37.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_38.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_38.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_38.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_38.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_39.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_39.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_39.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_39.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_4.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_4.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_4.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_40.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_40.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_40.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_40.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_41.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_41.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_41.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_41.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_42.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_42.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_42.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_42.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_43.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_43.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_43.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_43.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_44.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_44.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_44.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_44.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_45.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_45.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_45.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_45.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_46.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_46.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_46.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_46.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_47.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_47.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_47.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_47.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_48.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_48.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_48.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_48.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_49.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_49.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_49.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_49.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_5.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_5.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_5.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_50.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_50.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_50.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_50.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_51.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_51.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_51.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_51.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_52.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_52.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_52.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_52.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_53.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_53.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_53.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_53.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_54.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_54.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_54.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_54.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_6.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_6.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_6.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_6.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_7.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_7.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_7.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_7.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_8.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_8.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_8.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_8.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_9.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_9.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_9.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_9.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_filter_0.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_filter_0.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_filter_0.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_filter_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_miodio_0.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_miodio_0.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_miodio_0.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_miodio_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_mode_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_mode_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_mode_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_mode_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_filter_1.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_filter_1.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_filter_1.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_filter_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_miodio_1.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_miodio_1.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_miodio_1.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_miodio_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_mode_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_mode_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_mode_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_mode_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_filter_2.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_filter_2.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_filter_2.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_filter_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_miodio_2.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_miodio_2.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_miodio_2.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_miodio_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_mode_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_mode_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_mode_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_mode_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_filter_3.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_filter_3.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_filter_3.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_filter_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_miodio_3.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_miodio_3.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_miodio_3.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_miodio_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_mode_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_mode_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_mode_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_mode_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_filter_4.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_filter_4.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_filter_4.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_filter_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_miodio_4.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_miodio_4.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_miodio_4.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_miodio_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_mode_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_mode_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_mode_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_mode_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_filter_5.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_filter_5.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_filter_5.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_filter_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_miodio_5.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_miodio_5.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_miodio_5.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_miodio_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_mode_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_mode_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_mode_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_mode_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_filter_6.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_filter_6.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_filter_6.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_filter_6.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_miodio_6.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_miodio_6.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_miodio_6.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_miodio_6.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_mode_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_mode_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_mode_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_mode_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_filter_7.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_filter_7.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_filter_7.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_filter_7.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_miodio_7.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_miodio_7.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_miodio_7.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_miodio_7.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_mode_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_mode_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_mode_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_mode_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.astate_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.astate_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.filter_activity.stored_value_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.filter_activity.stored_value_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.filter_activity.stored_vector_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.filter_activity.stored_vector_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[0].u_filter.stored_value_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[0].u_filter.stored_value_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[0].u_filter.stored_vector_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[0].u_filter.stored_vector_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[1].u_filter.stored_value_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[1].u_filter.stored_value_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[1].u_filter.stored_vector_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[1].u_filter.stored_vector_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[2].u_filter.stored_value_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[2].u_filter.stored_value_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[2].u_filter.stored_vector_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[2].u_filter.stored_vector_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.u_cdc_suspend_req.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.u_cdc_suspend_req.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.u_cdc_suspend_req.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.u_cdc_suspend_req.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.beat_ctr_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.beat_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.phase_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.phase_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.common_sync_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.common_sync_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.u_common_sync1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.u_common_sync1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.u_common_sync1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.u_common_sync1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.intg_err_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_0_x_0.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_0_x_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_0_x_0.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_0_x_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_0_y_0.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_0_y_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_0_y_0.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_0_y_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_1_x_1.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_1_x_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_1_x_1.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_1_x_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_1_y_1.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_1_y_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_1_y_1.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_1_y_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_2_x_2.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_2_x_2.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_2_x_2.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_2_x_2.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_2_y_2.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_2_y_2.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_2_y_2.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_2_y_2.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_3_x_3.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_3_x_3.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_3_x_3.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_3_x_3.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_3_y_3.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_3_y_3.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_3_y_3.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_3_y_3.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_4_x_4.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_4_x_4.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_4_x_4.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_4_x_4.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_4_y_4.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_4_y_4.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_4_y_4.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_4_y_4.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_5_x_5.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_5_x_5.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_5_x_5.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_5_x_5.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_5_y_5.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_5_y_5.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_5_y_5.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_5_y_5.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_clk_div.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_clk_div.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_clk_div.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_clk_div.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_cntr_en.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_cntr_en.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_cntr_en.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_cntr_en.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_dc_resn.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_dc_resn.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_dc_resn.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_dc_resn.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_0_a_0.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_0_a_0.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_0_a_0.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_0_a_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_0_b_0.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_0_b_0.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_0_b_0.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_0_b_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_1_a_1.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_1_a_1.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_1_a_1.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_1_a_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_1_b_1.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_1_b_1.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_1_b_1.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_1_b_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_2_a_2.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_2_a_2.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_2_a_2.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_2_a_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_2_b_2.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_2_b_2.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_2_b_2.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_2_b_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_3_a_3.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_3_a_3.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_3_a_3.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_3_a_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_3_b_3.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_3_b_3.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_3_b_3.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_3_b_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_4_a_4.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_4_a_4.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_4_a_4.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_4_a_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_4_b_4.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_4_b_4.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_4_b_4.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_4_b_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_5_a_5.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_5_a_5.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_5_a_5.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_5_a_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_5_b_5.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_5_b_5.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_5_b_5.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_5_b_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_0.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_0.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_0.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_1.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_1.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_1.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_2.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_2.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_2.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_3.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_3.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_3.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_4.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_4.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_4.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_5.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_5.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_5.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_0.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_0.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_0.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_1.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_1.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_1.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_2.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_2.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_2.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_3.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_3.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_3.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_4.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_4.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_4.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_5.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_5.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_5.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_blink_en_0.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_blink_en_0.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_blink_en_0.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_blink_en_0.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_htbt_en_0.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_htbt_en_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_htbt_en_0.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_htbt_en_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_phase_delay_0.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_phase_delay_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_phase_delay_0.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_phase_delay_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_blink_en_1.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_blink_en_1.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_blink_en_1.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_blink_en_1.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_htbt_en_1.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_htbt_en_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_htbt_en_1.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_htbt_en_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_phase_delay_1.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_phase_delay_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_phase_delay_1.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_phase_delay_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_blink_en_2.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_blink_en_2.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_blink_en_2.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_blink_en_2.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_htbt_en_2.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_htbt_en_2.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_htbt_en_2.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_htbt_en_2.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_phase_delay_2.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_phase_delay_2.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_phase_delay_2.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_phase_delay_2.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_blink_en_3.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_blink_en_3.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_blink_en_3.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_blink_en_3.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_htbt_en_3.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_htbt_en_3.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_htbt_en_3.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_htbt_en_3.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_phase_delay_3.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_phase_delay_3.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_phase_delay_3.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_phase_delay_3.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_blink_en_4.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_blink_en_4.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_blink_en_4.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_blink_en_4.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_htbt_en_4.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_htbt_en_4.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_htbt_en_4.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_htbt_en_4.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_phase_delay_4.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_phase_delay_4.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_phase_delay_4.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_phase_delay_4.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_blink_en_5.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_blink_en_5.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_blink_en_5.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_blink_en_5.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_htbt_en_5.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_htbt_en_5.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_htbt_en_5.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_htbt_en_5.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_phase_delay_5.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_phase_delay_5.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_phase_delay_5.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_phase_delay_5.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_regen.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_regen.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_regen.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_regen.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ack_pwrdn_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ack_pwrdn_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ack_pwrdn_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ack_pwrdn_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ack_pwrup_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ack_pwrup_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ack_pwrup_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ack_pwrup_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ast_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ast_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ast_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ast_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ext_req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ext_req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ext_req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ext_req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_pwrup_chg_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_pwrup_chg_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_pwrup_chg_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_pwrup_chg_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_req_pwrdn_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_req_pwrdn_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_req_pwrdn_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_req_pwrdn_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_req_pwrup_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_req_pwrup_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_req_pwrup_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_req_pwrup_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_scdc_sync.dst_level_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_scdc_sync.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_scdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_scdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_scdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_scdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_scdc_sync.src_level  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_scdc_sync.src_level   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.dst_level_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.src_level  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.src_level   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_ext_req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_ext_req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_ext_req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_ext_req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.pwrup_cause_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.pwrup_cause_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.pwrup_cause_toggle_q2  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.pwrup_cause_toggle_q2   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_ast_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_ast_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_ast_q2    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_ast_q2 &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_core_clk_en_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_core_clk_en_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_io_clk_en_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_io_clk_en_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_main_pd_no    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_main_pd_no &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_reset_en_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_reset_en_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_usb_clk_en_active_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_usb_clk_en_active_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_usb_clk_en_lp_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_usb_clk_en_lp_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_wakeup_en_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_wakeup_en_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_flash_idle.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_flash_idle.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_flash_idle.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_flash_idle.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_otp.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_otp.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_otp.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_otp.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_rom_ctrl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_rom_ctrl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_rom_ctrl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_rom_ctrl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.ack_pwrup_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.ack_pwrup_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.ip_clk_en_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.ip_clk_en_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.low_power_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.low_power_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.req_pwrdn_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.req_pwrdn_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.reset_cause_q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.reset_cause_q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.reset_ongoing_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.reset_ongoing_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.rst_lc_req_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.rst_lc_req_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.rst_sys_req_q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.rst_sys_req_q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.state_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.state_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.strap_sampled  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.strap_sampled   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_fetch_en.u_prim_flop.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_fetch_en.u_prim_flop.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_reg_lc_init.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_reg_lc_init.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_reg_otp_init.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_reg_otp_init.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_slow_sync_lc_done.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_slow_sync_lc_done.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_slow_sync_lc_done.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_slow_sync_lc_done.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_sync_lc_done.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_sync_lc_done.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_sync_lc_done.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_sync_lc_done.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.ack_pwrdn_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.ack_pwrdn_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.cause_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.cause_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.cause_toggle_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.cause_toggle_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.core_clk_en_q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.core_clk_en_q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.io_clk_en_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.io_clk_en_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.pd_nq == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.pd_nq  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.pwr_clamp_env_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.pwr_clamp_env_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.pwr_clamp_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.pwr_clamp_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.req_pwrup_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.req_pwrup_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.state_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.state_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.usb_clk_en_q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.usb_clk_en_q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_wake_info.info == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_wake_info.info  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_wake_info.record_en    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_wake_info.record_en &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_wake_info.start_capture_q1 == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_wake_info.start_capture_q1  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.intr_wakeup.intr_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.intr_wakeup.intr_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.lowpwr_cfg_wen   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.lowpwr_cfg_wen    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_esc_rx.state_q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_esc_rx.state_q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_esc_rx.u_decode_esc.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_esc_rx.u_decode_esc.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_esc_rx.u_decode_esc.level_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_esc_rx.u_decode_esc.level_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_esc_rx.u_prim_generic_flop.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_esc_rx.u_prim_generic_flop.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_cfg_cdc_sync.q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_cfg_cdc_sync.q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_cfg_cdc_sync.qe  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_cfg_cdc_sync.qe   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_core_clk_en.q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_core_clk_en.q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_core_clk_en.qe   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_core_clk_en.qe    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_io_clk_en.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_io_clk_en.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_io_clk_en.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_io_clk_en.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_low_power_hint.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_low_power_hint.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_low_power_hint.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_low_power_hint.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_main_pd_n.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_main_pd_n.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_main_pd_n.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_main_pd_n.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_active.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_active.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_active.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_active.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_lp.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_lp.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_lp.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_lp.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_escalate_reset_status.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_escalate_reset_status.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_escalate_reset_status.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_escalate_reset_status.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_intr_enable.q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_intr_enable.q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_intr_enable.qe   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_intr_enable.qe    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_intr_state.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_intr_state.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_intr_state.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_intr_state.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_en_0.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_en_0.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_en_0.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_en_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_en_1.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_en_1.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_en_1.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_en_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_regwen.q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_regwen.q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_regwen.qe   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_status_val_0.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_status_val_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_status_val_0.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_status_val_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_status_val_1.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_status_val_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_status_val_1.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_status_val_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_info_capture_dis.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_info_capture_dis.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_info_capture_dis.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_info_capture_dis.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_0.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_0.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_0.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_1.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_1.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_1.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_2.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_2.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_2.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_3.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_3.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_3.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_4.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_4.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_4.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_0.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_0.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_1.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_1.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_2.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_2.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_2.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_2.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_3.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_3.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_3.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_3.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_4.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_4.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_4.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_4.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_regwen.q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_regwen.q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_regwen.qe  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_regwen.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.first_reset  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.first_reset   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.cnt  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.cnt   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_filter_n == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_filter_n  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.u_rst_flop.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.u_rst_flop.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[0].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[0].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[0].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[0].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[1].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[1].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[1].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[1].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[2].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[2].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[2].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[2].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[3].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[3].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[3].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[3].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[4].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[4].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[4].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[4].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[5].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[5].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[5].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[5].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[6].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[6].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[6].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[6].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_lc_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_lc_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_lc_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_lc_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_device.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_device.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_device.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_device.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_host0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_host0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_host0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_host0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_host1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_host1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_host1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_host1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys_aon.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys_aon.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys_aon.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys_aon.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_alert_info.slots_q == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_alert_info.slots_q  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io_div2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io_div2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io_div2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io_div2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_sys_aon.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_sys_aon.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_sys_aon.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_sys_aon.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_sys_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_sys_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_sys_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_sys_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_cpu_info.slots_q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_cpu_info.slots_q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_cpu_reset_synced.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_cpu_reset_synced.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_cpu_reset_synced.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_cpu_reset_synced.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_lc_src.gen_rst_pd_n[0].u_pd_rst.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_lc_src.gen_rst_pd_n[0].u_pd_rst.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_lc_src.u_aon_rst.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_lc_src.u_aon_rst.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_lc_src.u_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_lc_src.u_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_lc_src.u_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_lc_src.u_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_info_ctrl_en.q == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_info_ctrl_en.q  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_info_ctrl_en.qe    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_info_ctrl_en.qe &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_info_ctrl_index.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_info_ctrl_index.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_info_ctrl_index.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_info_ctrl_index.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_regwen.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_regwen.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_regwen.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_regwen.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_en.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_en.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_en.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_en.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_index.q    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_index.q &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_index.qe   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_index.qe    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_regwen.q == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_regwen.qe    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_hw_req.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_hw_req.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_hw_req.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_hw_req.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_low_power_exit.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_low_power_exit.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_low_power_exit.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_low_power_exit.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_ndm_reset.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_ndm_reset.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_ndm_reset.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_ndm_reset.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_por.q == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_por.q  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_por.qe    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_por.qe &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_0.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_0.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_0.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_0.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_1.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_1.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_1.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_1.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_2.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_2.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_2.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_2.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_3.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_3.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_3.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_3.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_4.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_4.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_4.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_4.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_5.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_5.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_5.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_5.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_6.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_6.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_6.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_6.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sys_src.gen_rst_pd_n[0].u_pd_rst.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sys_src.gen_rst_pd_n[0].u_pd_rst.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sys_src.u_aon_rst.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sys_src.u_aon_rst.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sys_src.u_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sys_src.u_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sys_src.u_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sys_src.u_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rv_timer.gen_harts[0].u_core.tick_count == top_level_upec.top_earlgrey_2.u_rv_timer.gen_harts[0].u_core.tick_count  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.gen_harts[0].u_intr_hw.intr_o  == top_level_upec.top_earlgrey_2.u_rv_timer.gen_harts[0].u_intr_hw.intr_o   &&
        top_level_upec.top_earlgrey_1.u_rv_timer.gen_harts[1].u_core.tick_count == top_level_upec.top_earlgrey_2.u_rv_timer.gen_harts[1].u_core.tick_count  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.gen_harts[1].u_intr_hw.intr_o  == top_level_upec.top_earlgrey_2.u_rv_timer.gen_harts[1].u_intr_hw.intr_o   &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_cfg0_prescale.q    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_cfg0_prescale.q &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_cfg0_prescale.qe   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_cfg0_prescale.qe    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_cfg0_step.q    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_cfg0_step.q &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_cfg0_step.qe   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_cfg0_step.qe    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_compare_lower0_0.q == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_compare_lower0_0.q  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_compare_lower0_0.qe    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_compare_lower0_0.qe &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_compare_upper0_0.q == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_compare_upper0_0.q  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_compare_upper0_0.qe    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_compare_upper0_0.qe &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_ctrl.q == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_ctrl.q  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_ctrl.qe    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_ctrl.qe &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_intr_enable0.q == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_intr_enable0.q  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_intr_enable0.qe    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_intr_enable0.qe &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_intr_state0.q  == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_intr_state0.q   &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_intr_state0.qe == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_intr_state0.qe  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_timer_v_lower0.q   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_timer_v_lower0.q    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_timer_v_lower0.qe  == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_timer_v_lower0.qe   &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_timer_v_upper0.q   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_timer_v_upper0.q    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_timer_v_upper0.qe  == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_timer_v_upper0.qe   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.intg_err_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_0.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_0.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_0.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_1.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_1.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_1.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_10.q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_10.q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_10.qe  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_10.qe   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_2.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_2.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_2.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_2.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_3.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_3.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_3.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_3.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_4.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_4.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_4.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_4.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_5.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_5.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_5.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_5.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_6.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_6.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_6.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_6.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_7.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_7.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_7.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_7.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_8.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_8.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_8.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_8.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_9.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_9.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_9.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_9.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_0.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_0.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_0.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_0.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_1.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_1.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_1.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_1.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_10.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_10.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_10.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_10.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_2.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_2.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_2.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_2.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_3.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_3.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_3.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_3.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_4.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_4.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_4.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_4.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_5.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_5.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_5.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_5.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_6.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_6.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_6.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_6.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_7.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_7.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_7.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_7.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_8.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_8.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_8.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_8.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_9.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_9.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_9.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_9.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_0.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_0.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_0.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_0.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_1.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_1.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_1.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_1.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_10.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_10.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_10.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_10.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_2.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_2.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_2.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_2.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_3.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_3.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_3.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_3.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_4.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_4.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_4.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_4.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_5.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_5.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_5.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_5.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_6.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_6.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_6.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_6.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_7.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_7.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_7.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_7.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_8.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_8.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_8.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_8.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_9.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_9.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_9.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_9.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_cfg_regwen.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_cfg_regwen.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_cfg_regwen.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_cfg_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_status_ast_init_done.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_status_ast_init_done.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_status_ast_init_done.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_status_ast_init_done.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_status_io_pok.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_status_io_pok.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_status_io_pok.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_status_io_pok.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.cmd_dp_sel_outclk    == top_level_upec.top_earlgrey_2.u_spi_device.cmd_dp_sel_outclk &&
        top_level_upec.top_earlgrey_1.u_spi_device.fwm_rxerr_q  == top_level_upec.top_earlgrey_2.u_spi_device.fwm_rxerr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.alert_set_q  == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.ping_set_q   == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.state_q  == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.state_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q    == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.io_mode_outclk   == top_level_upec.top_earlgrey_2.u_spi_device.io_mode_outclk    &&
        top_level_upec.top_earlgrey_1.u_spi_device.rxf_full_q   == top_level_upec.top_earlgrey_2.u_spi_device.rxf_full_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.rxlvl    == top_level_upec.top_earlgrey_2.u_spi_device.rxlvl &&
        top_level_upec.top_earlgrey_1.u_spi_device.sram_rxf_full_q  == top_level_upec.top_earlgrey_2.u_spi_device.sram_rxf_full_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.txf_empty_q  == top_level_upec.top_earlgrey_2.u_spi_device.txf_empty_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.txlvl    == top_level_upec.top_earlgrey_2.u_spi_device.txlvl &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_cmdparse.opcode_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_cmdparse.opcode_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_cmdparse.st    == top_level_upec.top_earlgrey_2.u_spi_device.u_cmdparse.st &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_fwmode_arb.gen_arb_ppc.u_reqarb.gen_normal_case.mask  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_fwmode_arb.gen_arb_ppc.u_reqarb.gen_normal_case.mask   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_gray_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_sync_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_sync_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.fifo_wptr_gray_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.fifo_wptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.fifo_wptr_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.fifo_wptr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.storage   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.byte_enable  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.byte_enable   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.cur_timer    == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.cur_timer &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.pos  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.pos   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.sram_req == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.sram_req  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.sram_wdata   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.sram_wdata    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.sram_write   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.sram_write    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.st   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.st    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.wptr == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.wptr  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_gray_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_sync_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_sync_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.fifo_wptr_gray_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.fifo_wptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.fifo_wptr_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.fifo_wptr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.storage   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.pos  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.pos   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.rptr == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.rptr  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.sram_rdata_q == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.sram_rdata_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.sram_req == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.sram_req  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.st   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.st    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.wptr_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.wptr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.a_rvalid_sram_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.a_rvalid_sram_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.b_rvalid_sram_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.b_rvalid_sram_q   &&
       // top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o   == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o    &&
       // top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o   == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o    &&
       // top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.mem == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.mem  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_p2s.cnt    == top_level_upec.top_earlgrey_2.u_spi_device.u_p2s.cnt &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_p2s.io_mode    == top_level_upec.top_earlgrey_2.u_spi_device.u_p2s.io_mode &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_p2s.out_shift  == top_level_upec.top_earlgrey_2.u_spi_device.u_p2s.out_shift   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_p2s.tx_state   == top_level_upec.top_earlgrey_2.u_spi_device.u_p2s.tx_state    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.addr_phase_outclk  == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.addr_phase_outclk   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.addrcnt    == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.addrcnt &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.addrcnt_outclk == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.addrcnt_outclk  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.bitcnt == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.bitcnt  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.cmd_filter == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.cmd_filter  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.cmd_info   == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.cmd_info    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.cmd_info_7th   == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.cmd_info_7th    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.csb_deassert   == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.csb_deassert    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.csb_deassert_outclk    == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.csb_deassert_outclk &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.dummycnt   == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.dummycnt    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.host_s_en_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.host_s_en_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.mailbox_hit    == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.mailbox_hit &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.opcode == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.opcode  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.passthrough_s_en   == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.passthrough_s_en    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.st == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.st  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.addr_q == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.addr_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.bitcnt == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.bitcnt  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.dummycnt   == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.dummycnt    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.fifo_byteoffset    == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.fifo_byteoffset &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.main_st    == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.main_st &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.p2s_byte_o == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.p2s_byte_o  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.p2s_valid_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.p2s_valid_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.readbuf_idx    == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.readbuf_idx &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_addr_swap_data.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_addr_swap_data.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_addr_swap_data.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_addr_swap_data.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_addr_swap_mask.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_addr_swap_mask.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_addr_swap_mask.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_addr_swap_mask.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_addr_4b_en.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_addr_4b_en.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_addr_4b_en.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_addr_4b_en.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_cpha.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_cpha.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_cpha.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_cpha.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_cpol.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_cpol.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_cpol.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_cpol.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_rx_order.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_rx_order.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_rx_order.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_rx_order.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_timer_v.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_timer_v.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_timer_v.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_timer_v.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_tx_order.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_tx_order.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_tx_order.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_tx_order.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_0.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_0.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_0.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_0.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_1.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_1.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_1.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_1.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_10.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_10.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_10.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_10.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_11.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_11.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_11.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_11.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_12.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_12.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_12.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_12.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_13.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_13.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_13.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_13.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_14.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_14.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_14.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_14.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_15.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_15.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_15.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_15.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_16.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_16.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_16.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_16.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_17.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_17.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_17.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_17.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_18.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_18.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_18.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_18.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_19.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_19.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_19.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_19.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_2.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_2.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_2.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_2.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_20.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_20.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_20.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_20.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_21.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_21.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_21.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_21.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_22.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_22.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_22.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_22.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_23.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_23.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_23.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_23.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_24.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_24.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_24.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_24.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_25.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_25.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_25.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_25.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_26.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_26.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_26.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_26.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_27.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_27.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_27.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_27.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_28.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_28.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_28.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_28.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_29.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_29.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_29.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_29.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_3.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_3.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_3.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_3.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_30.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_30.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_30.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_30.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_31.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_31.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_31.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_31.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_4.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_4.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_4.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_4.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_5.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_5.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_5.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_5.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_6.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_6.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_6.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_6.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_7.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_7.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_7.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_7.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_8.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_8.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_8.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_8.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_9.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_9.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_9.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_9.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_32.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_32.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_32.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_32.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_33.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_33.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_33.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_33.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_34.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_34.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_34.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_34.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_35.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_35.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_35.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_35.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_36.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_36.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_36.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_36.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_37.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_37.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_37.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_37.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_38.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_38.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_38.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_38.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_39.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_39.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_39.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_39.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_40.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_40.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_40.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_40.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_41.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_41.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_41.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_41.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_42.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_42.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_42.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_42.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_43.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_43.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_43.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_43.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_44.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_44.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_44.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_44.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_45.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_45.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_45.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_45.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_46.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_46.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_46.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_46.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_47.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_47.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_47.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_47.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_48.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_48.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_48.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_48.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_49.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_49.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_49.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_49.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_50.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_50.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_50.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_50.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_51.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_51.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_51.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_51.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_52.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_52.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_52.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_52.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_53.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_53.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_53.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_53.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_54.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_54.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_54.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_54.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_55.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_55.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_55.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_55.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_56.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_56.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_56.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_56.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_57.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_57.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_57.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_57.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_58.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_58.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_58.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_58.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_59.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_59.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_59.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_59.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_60.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_60.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_60.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_60.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_61.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_61.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_61.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_61.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_62.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_62.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_62.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_62.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_63.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_63.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_63.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_63.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_64.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_64.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_64.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_64.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_65.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_65.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_65.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_65.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_66.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_66.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_66.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_66.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_67.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_67.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_67.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_67.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_68.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_68.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_68.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_68.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_69.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_69.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_69.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_69.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_70.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_70.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_70.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_70.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_71.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_71.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_71.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_71.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_72.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_72.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_72.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_72.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_73.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_73.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_73.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_73.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_74.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_74.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_74.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_74.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_75.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_75.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_75.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_75.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_76.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_76.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_76.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_76.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_77.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_77.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_77.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_77.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_78.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_78.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_78.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_78.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_79.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_79.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_79.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_79.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_80.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_80.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_80.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_80.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_81.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_81.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_81.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_81.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_82.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_82.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_82.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_82.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_83.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_83.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_83.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_83.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_84.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_84.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_84.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_84.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_85.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_85.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_85.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_85.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_86.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_86.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_86.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_86.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_87.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_87.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_87.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_87.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_88.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_88.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_88.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_88.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_89.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_89.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_89.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_89.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_90.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_90.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_90.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_90.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_91.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_91.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_91.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_91.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_92.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_92.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_92.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_92.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_93.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_93.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_93.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_93.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_94.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_94.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_94.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_94.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_95.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_95.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_95.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_95.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_100.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_100.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_100.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_100.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_101.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_101.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_101.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_101.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_102.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_102.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_102.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_102.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_103.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_103.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_103.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_103.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_104.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_104.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_104.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_104.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_105.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_105.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_105.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_105.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_106.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_106.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_106.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_106.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_107.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_107.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_107.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_107.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_108.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_108.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_108.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_108.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_109.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_109.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_109.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_109.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_110.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_110.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_110.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_110.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_111.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_111.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_111.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_111.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_112.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_112.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_112.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_112.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_113.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_113.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_113.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_113.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_114.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_114.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_114.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_114.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_115.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_115.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_115.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_115.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_116.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_116.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_116.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_116.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_117.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_117.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_117.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_117.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_118.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_118.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_118.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_118.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_119.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_119.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_119.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_119.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_120.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_120.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_120.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_120.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_121.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_121.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_121.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_121.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_122.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_122.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_122.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_122.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_123.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_123.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_123.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_123.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_124.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_124.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_124.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_124.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_125.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_125.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_125.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_125.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_126.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_126.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_126.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_126.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_127.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_127.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_127.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_127.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_96.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_96.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_96.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_96.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_97.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_97.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_97.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_97.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_98.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_98.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_98.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_98.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_99.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_99.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_99.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_99.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_128.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_128.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_128.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_128.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_129.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_129.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_129.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_129.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_130.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_130.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_130.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_130.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_131.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_131.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_131.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_131.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_132.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_132.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_132.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_132.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_133.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_133.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_133.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_133.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_134.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_134.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_134.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_134.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_135.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_135.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_135.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_135.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_136.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_136.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_136.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_136.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_137.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_137.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_137.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_137.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_138.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_138.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_138.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_138.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_139.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_139.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_139.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_139.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_140.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_140.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_140.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_140.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_141.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_141.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_141.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_141.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_142.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_142.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_142.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_142.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_143.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_143.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_143.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_143.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_144.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_144.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_144.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_144.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_145.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_145.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_145.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_145.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_146.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_146.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_146.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_146.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_147.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_147.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_147.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_147.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_148.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_148.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_148.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_148.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_149.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_149.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_149.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_149.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_150.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_150.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_150.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_150.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_151.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_151.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_151.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_151.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_152.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_152.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_152.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_152.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_153.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_153.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_153.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_153.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_154.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_154.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_154.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_154.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_155.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_155.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_155.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_155.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_156.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_156.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_156.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_156.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_157.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_157.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_157.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_157.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_158.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_158.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_158.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_158.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_159.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_159.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_159.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_159.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_160.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_160.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_160.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_160.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_161.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_161.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_161.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_161.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_162.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_162.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_162.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_162.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_163.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_163.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_163.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_163.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_164.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_164.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_164.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_164.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_165.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_165.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_165.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_165.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_166.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_166.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_166.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_166.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_167.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_167.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_167.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_167.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_168.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_168.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_168.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_168.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_169.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_169.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_169.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_169.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_170.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_170.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_170.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_170.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_171.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_171.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_171.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_171.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_172.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_172.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_172.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_172.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_173.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_173.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_173.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_173.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_174.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_174.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_174.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_174.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_175.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_175.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_175.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_175.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_176.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_176.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_176.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_176.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_177.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_177.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_177.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_177.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_178.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_178.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_178.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_178.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_179.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_179.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_179.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_179.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_180.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_180.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_180.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_180.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_181.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_181.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_181.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_181.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_182.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_182.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_182.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_182.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_183.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_183.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_183.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_183.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_184.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_184.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_184.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_184.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_185.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_185.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_185.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_185.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_186.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_186.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_186.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_186.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_187.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_187.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_187.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_187.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_188.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_188.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_188.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_188.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_189.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_189.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_189.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_189.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_190.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_190.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_190.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_190.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_191.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_191.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_191.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_191.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_192.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_192.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_192.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_192.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_193.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_193.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_193.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_193.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_194.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_194.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_194.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_194.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_195.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_195.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_195.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_195.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_196.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_196.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_196.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_196.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_197.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_197.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_197.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_197.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_198.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_198.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_198.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_198.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_199.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_199.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_199.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_199.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_200.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_200.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_200.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_200.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_201.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_201.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_201.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_201.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_202.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_202.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_202.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_202.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_203.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_203.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_203.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_203.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_204.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_204.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_204.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_204.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_205.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_205.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_205.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_205.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_206.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_206.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_206.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_206.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_207.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_207.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_207.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_207.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_208.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_208.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_208.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_208.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_209.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_209.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_209.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_209.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_210.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_210.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_210.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_210.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_211.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_211.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_211.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_211.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_212.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_212.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_212.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_212.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_213.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_213.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_213.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_213.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_214.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_214.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_214.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_214.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_215.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_215.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_215.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_215.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_216.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_216.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_216.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_216.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_217.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_217.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_217.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_217.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_218.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_218.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_218.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_218.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_219.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_219.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_219.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_219.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_220.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_220.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_220.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_220.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_221.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_221.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_221.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_221.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_222.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_222.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_222.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_222.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_223.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_223.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_223.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_223.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_224.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_224.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_224.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_224.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_225.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_225.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_225.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_225.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_226.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_226.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_226.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_226.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_227.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_227.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_227.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_227.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_228.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_228.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_228.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_228.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_229.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_229.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_229.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_229.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_230.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_230.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_230.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_230.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_231.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_231.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_231.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_231.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_232.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_232.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_232.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_232.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_233.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_233.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_233.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_233.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_234.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_234.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_234.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_234.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_235.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_235.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_235.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_235.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_236.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_236.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_236.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_236.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_237.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_237.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_237.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_237.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_238.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_238.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_238.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_238.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_239.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_239.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_239.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_239.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_240.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_240.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_240.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_240.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_241.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_241.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_241.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_241.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_242.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_242.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_242.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_242.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_243.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_243.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_243.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_243.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_244.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_244.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_244.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_244.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_245.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_245.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_245.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_245.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_246.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_246.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_246.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_246.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_247.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_247.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_247.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_247.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_248.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_248.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_248.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_248.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_249.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_249.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_249.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_249.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_250.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_250.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_250.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_250.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_251.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_251.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_251.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_251.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_252.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_252.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_252.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_252.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_253.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_253.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_253.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_253.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_254.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_254.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_254.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_254.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_255.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_255.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_255.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_255.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_4b_affected_0.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_4b_affected_0.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_4b_affected_0.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_4b_affected_0.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_en_0.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_en_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_en_0.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_en_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_swap_en_0.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_swap_en_0.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_swap_en_0.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_swap_en_0.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_dummy_en_0.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_dummy_en_0.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_dummy_en_0.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_dummy_en_0.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_dummy_size_0.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_dummy_size_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_dummy_size_0.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_dummy_size_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_opcode_0.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_opcode_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_opcode_0.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_opcode_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_payload_dir_0.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_payload_dir_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_payload_dir_0.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_payload_dir_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_payload_en_0.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_payload_en_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_payload_en_0.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_payload_en_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_4b_affected_10.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_4b_affected_10.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_4b_affected_10.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_4b_affected_10.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_en_10.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_en_10.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_en_10.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_en_10.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_swap_en_10.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_swap_en_10.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_swap_en_10.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_swap_en_10.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_dummy_en_10.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_dummy_en_10.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_dummy_en_10.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_dummy_en_10.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_dummy_size_10.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_dummy_size_10.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_dummy_size_10.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_dummy_size_10.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_opcode_10.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_opcode_10.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_opcode_10.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_opcode_10.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_payload_dir_10.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_payload_dir_10.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_payload_dir_10.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_payload_dir_10.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_payload_en_10.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_payload_en_10.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_payload_en_10.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_payload_en_10.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_4b_affected_11.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_4b_affected_11.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_4b_affected_11.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_4b_affected_11.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_en_11.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_en_11.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_en_11.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_en_11.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_swap_en_11.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_swap_en_11.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_swap_en_11.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_swap_en_11.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_dummy_en_11.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_dummy_en_11.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_dummy_en_11.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_dummy_en_11.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_dummy_size_11.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_dummy_size_11.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_dummy_size_11.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_dummy_size_11.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_opcode_11.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_opcode_11.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_opcode_11.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_opcode_11.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_payload_dir_11.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_payload_dir_11.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_payload_dir_11.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_payload_dir_11.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_payload_en_11.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_payload_en_11.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_payload_en_11.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_payload_en_11.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_4b_affected_12.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_4b_affected_12.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_4b_affected_12.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_4b_affected_12.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_en_12.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_en_12.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_en_12.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_en_12.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_swap_en_12.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_swap_en_12.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_swap_en_12.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_swap_en_12.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_dummy_en_12.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_dummy_en_12.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_dummy_en_12.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_dummy_en_12.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_dummy_size_12.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_dummy_size_12.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_dummy_size_12.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_dummy_size_12.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_opcode_12.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_opcode_12.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_opcode_12.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_opcode_12.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_payload_dir_12.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_payload_dir_12.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_payload_dir_12.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_payload_dir_12.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_payload_en_12.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_payload_en_12.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_payload_en_12.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_payload_en_12.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_4b_affected_13.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_4b_affected_13.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_4b_affected_13.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_4b_affected_13.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_en_13.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_en_13.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_en_13.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_en_13.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_swap_en_13.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_swap_en_13.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_swap_en_13.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_swap_en_13.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_dummy_en_13.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_dummy_en_13.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_dummy_en_13.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_dummy_en_13.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_dummy_size_13.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_dummy_size_13.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_dummy_size_13.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_dummy_size_13.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_opcode_13.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_opcode_13.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_opcode_13.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_opcode_13.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_payload_dir_13.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_payload_dir_13.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_payload_dir_13.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_payload_dir_13.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_payload_en_13.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_payload_en_13.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_payload_en_13.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_payload_en_13.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_4b_affected_14.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_4b_affected_14.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_4b_affected_14.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_4b_affected_14.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_en_14.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_en_14.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_en_14.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_en_14.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_swap_en_14.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_swap_en_14.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_swap_en_14.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_swap_en_14.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_dummy_en_14.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_dummy_en_14.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_dummy_en_14.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_dummy_en_14.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_dummy_size_14.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_dummy_size_14.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_dummy_size_14.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_dummy_size_14.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_opcode_14.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_opcode_14.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_opcode_14.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_opcode_14.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_payload_dir_14.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_payload_dir_14.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_payload_dir_14.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_payload_dir_14.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_payload_en_14.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_payload_en_14.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_payload_en_14.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_payload_en_14.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_4b_affected_15.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_4b_affected_15.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_4b_affected_15.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_4b_affected_15.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_en_15.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_en_15.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_en_15.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_en_15.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_swap_en_15.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_swap_en_15.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_swap_en_15.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_swap_en_15.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_dummy_en_15.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_dummy_en_15.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_dummy_en_15.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_dummy_en_15.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_dummy_size_15.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_dummy_size_15.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_dummy_size_15.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_dummy_size_15.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_opcode_15.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_opcode_15.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_opcode_15.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_opcode_15.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_payload_dir_15.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_payload_dir_15.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_payload_dir_15.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_payload_dir_15.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_payload_en_15.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_payload_en_15.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_payload_en_15.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_payload_en_15.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_4b_affected_1.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_4b_affected_1.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_4b_affected_1.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_4b_affected_1.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_en_1.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_en_1.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_en_1.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_en_1.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_swap_en_1.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_swap_en_1.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_swap_en_1.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_swap_en_1.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_dummy_en_1.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_dummy_en_1.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_dummy_en_1.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_dummy_en_1.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_dummy_size_1.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_dummy_size_1.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_dummy_size_1.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_dummy_size_1.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_opcode_1.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_opcode_1.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_opcode_1.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_opcode_1.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_payload_dir_1.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_payload_dir_1.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_payload_dir_1.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_payload_dir_1.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_payload_en_1.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_payload_en_1.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_payload_en_1.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_payload_en_1.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_4b_affected_2.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_4b_affected_2.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_4b_affected_2.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_4b_affected_2.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_en_2.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_en_2.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_en_2.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_en_2.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_swap_en_2.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_swap_en_2.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_swap_en_2.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_swap_en_2.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_dummy_en_2.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_dummy_en_2.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_dummy_en_2.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_dummy_en_2.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_dummy_size_2.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_dummy_size_2.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_dummy_size_2.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_dummy_size_2.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_opcode_2.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_opcode_2.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_opcode_2.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_opcode_2.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_payload_dir_2.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_payload_dir_2.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_payload_dir_2.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_payload_dir_2.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_payload_en_2.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_payload_en_2.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_payload_en_2.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_payload_en_2.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_4b_affected_3.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_4b_affected_3.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_4b_affected_3.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_4b_affected_3.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_en_3.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_en_3.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_en_3.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_en_3.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_swap_en_3.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_swap_en_3.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_swap_en_3.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_swap_en_3.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_dummy_en_3.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_dummy_en_3.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_dummy_en_3.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_dummy_en_3.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_dummy_size_3.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_dummy_size_3.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_dummy_size_3.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_dummy_size_3.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_opcode_3.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_opcode_3.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_opcode_3.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_opcode_3.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_payload_dir_3.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_payload_dir_3.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_payload_dir_3.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_payload_dir_3.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_payload_en_3.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_payload_en_3.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_payload_en_3.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_payload_en_3.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_4b_affected_4.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_4b_affected_4.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_4b_affected_4.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_4b_affected_4.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_en_4.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_en_4.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_en_4.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_en_4.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_swap_en_4.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_swap_en_4.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_swap_en_4.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_swap_en_4.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_dummy_en_4.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_dummy_en_4.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_dummy_en_4.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_dummy_en_4.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_dummy_size_4.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_dummy_size_4.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_dummy_size_4.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_dummy_size_4.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_opcode_4.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_opcode_4.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_opcode_4.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_opcode_4.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_payload_dir_4.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_payload_dir_4.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_payload_dir_4.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_payload_dir_4.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_payload_en_4.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_payload_en_4.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_payload_en_4.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_payload_en_4.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_4b_affected_5.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_4b_affected_5.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_4b_affected_5.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_4b_affected_5.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_en_5.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_en_5.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_en_5.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_en_5.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_swap_en_5.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_swap_en_5.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_swap_en_5.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_swap_en_5.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_dummy_en_5.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_dummy_en_5.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_dummy_en_5.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_dummy_en_5.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_dummy_size_5.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_dummy_size_5.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_dummy_size_5.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_dummy_size_5.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_opcode_5.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_opcode_5.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_opcode_5.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_opcode_5.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_payload_dir_5.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_payload_dir_5.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_payload_dir_5.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_payload_dir_5.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_payload_en_5.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_payload_en_5.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_payload_en_5.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_payload_en_5.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_4b_affected_6.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_4b_affected_6.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_4b_affected_6.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_4b_affected_6.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_en_6.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_en_6.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_en_6.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_en_6.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_swap_en_6.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_swap_en_6.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_swap_en_6.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_swap_en_6.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_dummy_en_6.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_dummy_en_6.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_dummy_en_6.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_dummy_en_6.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_dummy_size_6.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_dummy_size_6.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_dummy_size_6.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_dummy_size_6.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_opcode_6.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_opcode_6.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_opcode_6.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_opcode_6.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_payload_dir_6.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_payload_dir_6.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_payload_dir_6.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_payload_dir_6.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_payload_en_6.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_payload_en_6.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_payload_en_6.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_payload_en_6.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_4b_affected_7.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_4b_affected_7.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_4b_affected_7.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_4b_affected_7.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_en_7.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_en_7.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_en_7.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_en_7.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_swap_en_7.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_swap_en_7.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_swap_en_7.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_swap_en_7.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_dummy_en_7.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_dummy_en_7.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_dummy_en_7.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_dummy_en_7.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_dummy_size_7.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_dummy_size_7.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_dummy_size_7.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_dummy_size_7.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_opcode_7.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_opcode_7.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_opcode_7.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_opcode_7.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_payload_dir_7.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_payload_dir_7.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_payload_dir_7.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_payload_dir_7.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_payload_en_7.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_payload_en_7.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_payload_en_7.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_payload_en_7.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_4b_affected_8.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_4b_affected_8.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_4b_affected_8.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_4b_affected_8.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_en_8.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_en_8.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_en_8.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_en_8.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_swap_en_8.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_swap_en_8.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_swap_en_8.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_swap_en_8.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_dummy_en_8.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_dummy_en_8.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_dummy_en_8.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_dummy_en_8.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_dummy_size_8.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_dummy_size_8.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_dummy_size_8.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_dummy_size_8.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_opcode_8.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_opcode_8.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_opcode_8.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_opcode_8.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_payload_dir_8.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_payload_dir_8.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_payload_dir_8.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_payload_dir_8.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_payload_en_8.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_payload_en_8.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_payload_en_8.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_payload_en_8.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_4b_affected_9.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_4b_affected_9.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_4b_affected_9.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_4b_affected_9.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_en_9.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_en_9.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_en_9.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_en_9.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_swap_en_9.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_swap_en_9.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_swap_en_9.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_swap_en_9.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_dummy_en_9.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_dummy_en_9.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_dummy_en_9.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_dummy_en_9.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_dummy_size_9.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_dummy_size_9.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_dummy_size_9.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_dummy_size_9.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_opcode_9.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_opcode_9.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_opcode_9.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_opcode_9.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_payload_dir_9.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_payload_dir_9.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_payload_dir_9.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_payload_dir_9.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_payload_en_9.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_payload_en_9.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_payload_en_9.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_payload_en_9.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_abort.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_abort.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_abort.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_abort.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_mode.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_mode.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_mode.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_mode.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_rst_rxfifo.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_rst_rxfifo.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_rst_rxfifo.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_rst_rxfifo.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_rst_txfifo.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_rst_txfifo.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_rst_txfifo.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_rst_txfifo.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_sram_clk_en.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_sram_clk_en.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_sram_clk_en.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_sram_clk_en.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_fifo_level_rxlvl.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_fifo_level_rxlvl.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_fifo_level_rxlvl.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_fifo_level_rxlvl.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_fifo_level_txlvl.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_fifo_level_txlvl.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_fifo_level_txlvl.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_fifo_level_txlvl.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxerr.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxerr.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxerr.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxerr.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxf.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxf.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxf.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxf.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxlvl.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxlvl.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxlvl.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxlvl.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxoverflow.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxoverflow.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxoverflow.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxoverflow.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_txlvl.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_txlvl.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_txlvl.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_txlvl.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_txunderflow.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_txunderflow.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_txunderflow.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_txunderflow.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxerr.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxerr.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxerr.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxerr.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxf.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxf.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxf.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxf.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxlvl.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxlvl.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxlvl.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxlvl.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxoverflow.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxoverflow.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxoverflow.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxoverflow.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_txlvl.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_txlvl.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_txlvl.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_txlvl.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_txunderflow.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_txunderflow.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_txunderflow.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_txunderflow.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_addr_base.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_addr_base.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_addr_base.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_addr_base.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_addr_limit.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_addr_limit.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_addr_limit.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_addr_limit.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_ptr_rptr.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_ptr_rptr.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_ptr_rptr.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_ptr_rptr.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_ptr_wptr.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_ptr_wptr.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_ptr_wptr.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_ptr_wptr.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.dev_select_outstanding    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.dev_select_outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.err_resp.err_opcode   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.err_resp.err_opcode    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.err_resp.err_req_pending  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.err_resp.err_req_pending   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.err_resp.err_rsp_pending  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.err_resp.err_rsp_pending   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.err_resp.err_size == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.err_resp.err_size  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.err_resp.err_source   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.err_resp.err_source    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.num_req_outstanding   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.num_req_outstanding    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_addr_base.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_addr_base.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_addr_base.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_addr_base.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_addr_limit.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_addr_limit.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_addr_limit.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_addr_limit.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_ptr_rptr.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_ptr_rptr.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_ptr_rptr.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_ptr_rptr.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_ptr_wptr.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_ptr_wptr.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_ptr_wptr.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_ptr_wptr.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_rxf_overflow.dst_level_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_rxf_overflow.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_rxf_overflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_rxf_overflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_rxf_overflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_rxf_overflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_rxf_overflow.src_level == top_level_upec.top_earlgrey_2.u_spi_device.u_rxf_overflow.src_level  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_s2p.bitcnt == top_level_upec.top_earlgrey_2.u_spi_device.u_s2p.bitcnt  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_s2p.cnt    == top_level_upec.top_earlgrey_2.u_spi_device.u_s2p.cnt &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_s2p.data_q == top_level_upec.top_earlgrey_2.u_spi_device.u_s2p.data_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sram_clk_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_spi_device.u_sram_clk_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_csb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_csb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_csb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_csb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_rxf.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_rxf.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_rxf.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_rxf.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_txe.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_txe.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_txe.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_txe.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.intg_error_q == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.intg_error_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_txf_underflow.dst_level_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_txf_underflow.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_txf_underflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_device.u_txf_underflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_txf_underflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_device.u_txf_underflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_txf_underflow.src_level    == top_level_upec.top_earlgrey_2.u_spi_device.u_txf_underflow.src_level &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.idle_q    == top_level_upec.top_earlgrey_2.u_spi_host0.idle_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.intr_hw_error.intr_o  == top_level_upec.top_earlgrey_2.u_spi_host0.intr_hw_error.intr_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.intr_hw_spi_event.intr_o  == top_level_upec.top_earlgrey_2.u_spi_host0.intr_hw_spi_event.intr_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.ready_q   == top_level_upec.top_earlgrey_2.u_spi_host0.ready_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.rx_full_q == top_level_upec.top_earlgrey_2.u_spi_host0.rx_full_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.rx_wm_q   == top_level_upec.top_earlgrey_2.u_spi_host0.rx_wm_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.tx_empty_q    == top_level_upec.top_earlgrey_2.u_spi_host0.tx_empty_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.tx_wm_q   == top_level_upec.top_earlgrey_2.u_spi_host0.tx_wm_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.cdc_req_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.cdc_req_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.command_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.command_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_ack_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_ack_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_fsm_cs == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_fsm_cs == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_req_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_req_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_csaat.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_csaat.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_csaat.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_csaat.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_direction.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_direction.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_direction.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_direction.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_len.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_len.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_len.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_len.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_speed.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_speed.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_speed.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_speed.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_clkdiv_0.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_clkdiv_0.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_clkdiv_0.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_clkdiv_0.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_cpha_0.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_cpha_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_cpha_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_cpha_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_cpol_0.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_cpol_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_cpol_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_cpol_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csnidle_0.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csnidle_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csnidle_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csnidle_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csnlead_0.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csnlead_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csnlead_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csnlead_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csntrail_0.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csntrail_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csntrail_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csntrail_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_fullcyc_0.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_fullcyc_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_fullcyc_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_fullcyc_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_passthru.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_passthru.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_passthru.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_passthru.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_spien.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_spien.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_spien.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_spien.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_sw_rst.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_sw_rst.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_sw_rst.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_sw_rst.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_csid.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_csid.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_csid.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_csid.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_cmdbusy.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_cmdbusy.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_cmdbusy.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_cmdbusy.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_cmdinval.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_cmdinval.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_cmdinval.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_cmdinval.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_csidinval.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_csidinval.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_csidinval.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_csidinval.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_overflow.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_overflow.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_underflow.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_underflow.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_underflow.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_underflow.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_cmdbusy.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_cmdbusy.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_cmdbusy.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_cmdbusy.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_cmdinval.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_cmdinval.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_cmdinval.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_cmdinval.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_csidinval.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_csidinval.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_csidinval.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_csidinval.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_overflow.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_overflow.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_underflow.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_underflow.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_underflow.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_underflow.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_idle.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_idle.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_idle.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_idle.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_ready.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_ready.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_ready.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_ready.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_rxfull.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_rxfull.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_rxfull.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_rxfull.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_rxwm.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_rxwm.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_rxwm.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_rxwm.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_txempty.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_txempty.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_txempty.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_txempty.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_txwm.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_txwm.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_txwm.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_txwm.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_enable_error.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_enable_error.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_enable_error.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_enable_error.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_enable_spi_event.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_enable_spi_event.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_enable_spi_event.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_enable_spi_event.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_state_error.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_state_error.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_state_error.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_state_error.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_state_spi_event.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_state_spi_event.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_state_spi_event.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_state_spi_event.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.dev_select_outstanding == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.dev_select_outstanding  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.err_resp.err_opcode    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.err_resp.err_opcode &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.err_resp.err_req_pending   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.err_resp.err_req_pending    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.err_resp.err_rsp_pending   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.err_resp.err_rsp_pending    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.err_resp.err_size  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.err_resp.err_size   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.err_resp.err_source    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.err_resp.err_source &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.num_req_outstanding    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.num_req_outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_active.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_active.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_active.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_active.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_byteorder.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_byteorder.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_byteorder.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_byteorder.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_ready.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_ready.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_ready.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_ready.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxempty.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxempty.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxempty.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxempty.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxfull.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxfull.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxfull.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxfull.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxqd.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxqd.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxqd.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxqd.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxstall.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxstall.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxstall.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxstall.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxwm.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxwm.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxwm.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxwm.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txempty.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txempty.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txempty.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txempty.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txfull.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txfull.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txfull.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txfull.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txqd.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txqd.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txqd.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txqd.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txstall.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txstall.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txstall.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txstall.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txwm.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txwm.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txwm.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txwm.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.bit_cntr_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.bit_cntr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.bit_shifting_cpha1   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.bit_shifting_cpha1    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.byte_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.byte_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.byte_ending_cpha1    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.byte_ending_cpha1 &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.byte_starting_cpha1  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.byte_starting_cpha1   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.clk_cntr_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.clk_cntr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.clkdiv_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.clkdiv_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.cmd_rd_en_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.cmd_rd_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.cmd_speed_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.cmd_speed_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.cmd_wr_en_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.cmd_wr_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.cpha_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.cpha_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.cpol_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.cpol_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csaat_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csaat_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csb_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csb_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csid_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csid_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csnidle_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csnidle_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csnlead_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csnlead_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csntrail_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csntrail_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.full_cyc_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.full_cyc_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.idle_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.idle_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.lead_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.lead_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.sample_en_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.sample_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.sample_en_q2 == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.sample_en_q2  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.sck_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.sck_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.spi_host_st_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.spi_host_st_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.trail_cntr_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.trail_cntr_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_merge.last_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_merge.last_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_merge.u_packer.clr_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_merge.u_packer.clr_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_merge.u_packer.data_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_merge.u_packer.data_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_merge.u_packer.depth_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_merge.u_packer.depth_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_select.u_packer.clr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_select.u_packer.clr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_select.u_packer.data_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_select.u_packer.data_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_select.u_packer.depth_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_select.u_packer.depth_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_select.u_packer.gen_unpack_mode.ptr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_select.u_packer.gen_unpack_mode.ptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_shift_reg.rx_buf_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_shift_reg.rx_buf_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_shift_reg.rx_buf_valid_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_shift_reg.rx_buf_valid_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_shift_reg.sd_i_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_shift_reg.sd_i_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_shift_reg.sr_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_shift_reg.sr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host0.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host0.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host0.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host0.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.error  == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.error   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.outstanding    == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.rdata  == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.rdata   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.reqid  == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.reqid   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.reqsz  == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.reqsz   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.rspop  == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.rspop   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.idle_q    == top_level_upec.top_earlgrey_2.u_spi_host1.idle_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.intr_hw_error.intr_o  == top_level_upec.top_earlgrey_2.u_spi_host1.intr_hw_error.intr_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.intr_hw_spi_event.intr_o  == top_level_upec.top_earlgrey_2.u_spi_host1.intr_hw_spi_event.intr_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.ready_q   == top_level_upec.top_earlgrey_2.u_spi_host1.ready_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.rx_full_q == top_level_upec.top_earlgrey_2.u_spi_host1.rx_full_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.rx_wm_q   == top_level_upec.top_earlgrey_2.u_spi_host1.rx_wm_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.tx_empty_q    == top_level_upec.top_earlgrey_2.u_spi_host1.tx_empty_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.tx_wm_q   == top_level_upec.top_earlgrey_2.u_spi_host1.tx_wm_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.cdc_req_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.cdc_req_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.command_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.command_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_ack_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_ack_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_fsm_cs == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_fsm_cs == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_req_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_req_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_csaat.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_csaat.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_csaat.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_csaat.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_direction.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_direction.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_direction.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_direction.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_len.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_len.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_len.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_len.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_speed.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_speed.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_speed.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_speed.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_clkdiv_0.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_clkdiv_0.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_clkdiv_0.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_clkdiv_0.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_cpha_0.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_cpha_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_cpha_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_cpha_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_cpol_0.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_cpol_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_cpol_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_cpol_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csnidle_0.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csnidle_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csnidle_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csnidle_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csnlead_0.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csnlead_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csnlead_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csnlead_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csntrail_0.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csntrail_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csntrail_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csntrail_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_fullcyc_0.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_fullcyc_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_fullcyc_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_fullcyc_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_passthru.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_passthru.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_passthru.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_passthru.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_spien.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_spien.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_spien.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_spien.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_sw_rst.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_sw_rst.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_sw_rst.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_sw_rst.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_csid.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_csid.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_csid.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_csid.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_cmdbusy.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_cmdbusy.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_cmdbusy.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_cmdbusy.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_cmdinval.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_cmdinval.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_cmdinval.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_cmdinval.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_csidinval.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_csidinval.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_csidinval.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_csidinval.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_overflow.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_overflow.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_underflow.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_underflow.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_underflow.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_underflow.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_cmdbusy.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_cmdbusy.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_cmdbusy.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_cmdbusy.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_cmdinval.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_cmdinval.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_cmdinval.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_cmdinval.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_csidinval.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_csidinval.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_csidinval.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_csidinval.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_overflow.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_overflow.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_underflow.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_underflow.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_underflow.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_underflow.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_idle.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_idle.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_idle.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_idle.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_ready.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_ready.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_ready.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_ready.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_rxfull.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_rxfull.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_rxfull.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_rxfull.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_rxwm.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_rxwm.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_rxwm.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_rxwm.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_txempty.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_txempty.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_txempty.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_txempty.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_txwm.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_txwm.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_txwm.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_txwm.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_enable_error.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_enable_error.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_enable_error.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_enable_error.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_enable_spi_event.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_enable_spi_event.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_enable_spi_event.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_enable_spi_event.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_state_error.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_state_error.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_state_error.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_state_error.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_state_spi_event.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_state_spi_event.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_state_spi_event.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_state_spi_event.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.dev_select_outstanding == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.dev_select_outstanding  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.err_resp.err_opcode    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.err_resp.err_opcode &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.err_resp.err_req_pending   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.err_resp.err_req_pending    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.err_resp.err_rsp_pending   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.err_resp.err_rsp_pending    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.err_resp.err_size  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.err_resp.err_size   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.err_resp.err_source    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.err_resp.err_source &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.num_req_outstanding    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.num_req_outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_active.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_active.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_active.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_active.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_byteorder.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_byteorder.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_byteorder.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_byteorder.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_ready.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_ready.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_ready.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_ready.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxempty.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxempty.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxempty.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxempty.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxfull.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxfull.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxfull.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxfull.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxqd.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxqd.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxqd.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxqd.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxstall.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxstall.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxstall.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxstall.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxwm.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxwm.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxwm.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxwm.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txempty.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txempty.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txempty.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txempty.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txfull.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txfull.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txfull.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txfull.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txqd.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txqd.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txqd.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txqd.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txstall.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txstall.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txstall.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txstall.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txwm.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txwm.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txwm.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txwm.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.bit_cntr_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.bit_cntr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.bit_shifting_cpha1   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.bit_shifting_cpha1    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.byte_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.byte_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.byte_ending_cpha1    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.byte_ending_cpha1 &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.byte_starting_cpha1  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.byte_starting_cpha1   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.clk_cntr_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.clk_cntr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.clkdiv_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.clkdiv_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.cmd_rd_en_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.cmd_rd_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.cmd_speed_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.cmd_speed_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.cmd_wr_en_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.cmd_wr_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.cpha_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.cpha_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.cpol_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.cpol_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csaat_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csaat_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csb_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csb_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csid_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csid_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csnidle_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csnidle_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csnlead_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csnlead_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csntrail_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csntrail_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.full_cyc_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.full_cyc_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.idle_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.idle_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.lead_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.lead_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.sample_en_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.sample_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.sample_en_q2 == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.sample_en_q2  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.sck_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.sck_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.spi_host_st_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.spi_host_st_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.trail_cntr_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.trail_cntr_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_merge.last_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_merge.last_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_merge.u_packer.clr_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_merge.u_packer.clr_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_merge.u_packer.data_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_merge.u_packer.data_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_merge.u_packer.depth_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_merge.u_packer.depth_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_select.u_packer.clr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_select.u_packer.clr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_select.u_packer.data_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_select.u_packer.data_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_select.u_packer.depth_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_select.u_packer.depth_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_select.u_packer.gen_unpack_mode.ptr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_select.u_packer.gen_unpack_mode.ptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_shift_reg.rx_buf_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_shift_reg.rx_buf_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_shift_reg.rx_buf_valid_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_shift_reg.rx_buf_valid_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_shift_reg.sd_i_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_shift_reg.sd_i_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_shift_reg.sr_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_shift_reg.sr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host1.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host1.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host1.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host1.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.error  == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.error   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.outstanding    == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.rdata  == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.rdata   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.reqid  == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.reqid   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.reqsz  == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.reqsz   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.rspop  == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.rspop   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.escalated_q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.escalated_q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.alert_set_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.alert_set_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.alert_test_set_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.alert_test_set_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.ping_set_q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.ping_set_q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.state_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.state_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.level_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.level_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.level_q    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.level_q &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_prim_generic_flop.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_prim_generic_flop.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.alert_set_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.alert_set_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.alert_test_set_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.alert_test_set_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.ping_set_q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.ping_set_q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.state_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.state_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.level_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.level_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.level_q    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.level_q &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_prim_generic_flop.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_prim_generic_flop.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.init_q    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.init_q &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.key_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.key_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.key_req_pending_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.key_req_pending_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.key_seed_valid_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.key_seed_valid_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.key_valid_q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.key_valid_q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.nonce_q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.nonce_q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.parity_error_q    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.parity_error_q &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_ctrl_regwen.q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_ctrl_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_ctrl_regwen.qe    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_ctrl_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_error_address.q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_error_address.q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_error_address.qe  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_error_address.qe   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_exec.q    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_exec.q &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_exec.qe   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_exec.qe    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_exec_regwen.q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_exec_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_exec_regwen.qe    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_exec_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.cfg_auto_block_timer    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.cfg_auto_block_timer &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_en.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_en.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_en.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_en.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_gray_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_sync_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_sync_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_wptr_gray_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_wptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_wptr_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_wptr_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.storage  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.storage   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_pwrb_in_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_pwrb_in_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_pwrb_in_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_pwrb_in_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.cfg_combo_timer == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.cfg_combo_timer  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.cfg_debounce_timer  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.cfg_debounce_timer   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.storage    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.storage &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.storage    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.storage &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.storage    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.storage &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.storage    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.storage &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.bat_disable_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.bat_disable_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.cfg_ec_rst_timer   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.cfg_ec_rst_timer    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.combo_det_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.combo_det_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.ec_rst_l_int   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.ec_rst_l_int    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.ec_rst_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.ec_rst_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.gsc_rst_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.gsc_rst_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.storage == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.storage  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.bat_disable_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.bat_disable_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.cfg_ec_rst_timer   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.cfg_ec_rst_timer    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.combo_det_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.combo_det_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.ec_rst_l_int   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.ec_rst_l_int    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.ec_rst_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.ec_rst_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.gsc_rst_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.gsc_rst_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.storage == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.storage  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.bat_disable_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.bat_disable_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.cfg_ec_rst_timer   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.cfg_ec_rst_timer    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.combo_det_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.combo_det_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.ec_rst_l_int   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.ec_rst_l_int    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.ec_rst_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.ec_rst_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.gsc_rst_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.gsc_rst_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.storage == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.storage  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.bat_disable_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.bat_disable_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.cfg_ec_rst_timer   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.cfg_ec_rst_timer    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.combo_det_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.combo_det_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.ec_rst_l_int   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.ec_rst_l_int    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.ec_rst_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.ec_rst_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.gsc_rst_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.gsc_rst_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.storage == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.storage  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer1_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer1_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer2_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer2_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer_state_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer_state_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.trigger_h_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.trigger_h_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.trigger_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.trigger_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer1_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer1_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer2_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer2_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer_state_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer_state_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.trigger_h_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.trigger_h_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.trigger_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.trigger_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer1_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer1_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer2_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer2_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer_state_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer_state_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.trigger_h_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.trigger_h_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.trigger_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.trigger_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer1_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer1_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer2_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer2_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer_state_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer_state_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.trigger_h_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.trigger_h_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.trigger_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.trigger_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.storage    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.storage &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.dst_level_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.src_level == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.src_level  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.dst_level_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.src_level == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.src_level  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.dst_level_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.src_level == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.src_level  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.dst_level_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.src_level == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.src_level  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key0_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key0_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key0_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key0_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key1_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key1_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key1_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key1_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key2_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key2_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key2_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key2_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_intr.i_sysrst_ctrl_intr_o.intr_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_intr.i_sysrst_ctrl_intr_o.intr_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_ac_present_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_ac_present_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_ac_present_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_ac_present_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_bat_disable_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_bat_disable_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_bat_disable_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_bat_disable_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.ac_present_intr_h2l_det_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.ac_present_intr_h2l_det_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.ac_present_intr_l2h_det_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.ac_present_intr_l2h_det_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.cfg_key_intr_timer    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.cfg_key_intr_timer &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.ec_rst_l_intr_h2l_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.ec_rst_l_intr_h2l_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.ec_rst_l_intr_l2h_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.ec_rst_l_intr_l2h_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.dst_level_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.src_level    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.src_level &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.dst_level_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.src_level    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.src_level &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.timer_cnt_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.timer_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.timer_state_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.timer_state_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.trigger_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.trigger_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_gray_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_sync_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_sync_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_wptr_gray_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_wptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_wptr_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_wptr_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.storage  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.storage   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.dst_level_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.src_level  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.src_level   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.dst_level_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.src_level  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.src_level   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.dst_level_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.src_level  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.src_level   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.dst_level_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.src_level  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.src_level   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key0_intr_h2l_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key0_intr_h2l_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key0_intr_l2h_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key0_intr_l2h_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key1_intr_h2l_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key1_intr_h2l_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key1_intr_l2h_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key1_intr_l2h_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key2_intr_h2l_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key2_intr_h2l_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key2_intr_l2h_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key2_intr_l2h_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.pwrb_intr_h2l_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.pwrb_intr_h2l_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.pwrb_intr_l2h_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.pwrb_intr_l2h_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ac_present_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ac_present_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ac_present_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ac_present_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.intg_err_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_auto_block_enable.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_auto_block_enable.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_auto_block_enable.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_auto_block_enable.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_debounce_timer.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_debounce_timer.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_debounce_timer.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_debounce_timer.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_sel.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_sel.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_sel.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_sel.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_value.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_value.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_value.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_value.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_sel.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_sel.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_sel.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_sel.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_value.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_value.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_value.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_value.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_sel.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_sel.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_sel.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_sel.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_value.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_value.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_value.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_value.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_0.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_0.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_0.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_0.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_1.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_1.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_1.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_1.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_2.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_2.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_2.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_2.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_3.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_3.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_3.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_3.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_bat_disable_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_bat_disable_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_bat_disable_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_bat_disable_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_ec_rst_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_ec_rst_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_ec_rst_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_ec_rst_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_gsc_rst_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_gsc_rst_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_gsc_rst_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_gsc_rst_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_interrupt_0.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_interrupt_0.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_interrupt_0.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_interrupt_0.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_bat_disable_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_bat_disable_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_bat_disable_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_bat_disable_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_ec_rst_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_ec_rst_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_ec_rst_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_ec_rst_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_gsc_rst_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_gsc_rst_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_gsc_rst_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_gsc_rst_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_interrupt_1.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_interrupt_1.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_interrupt_1.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_interrupt_1.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_bat_disable_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_bat_disable_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_bat_disable_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_bat_disable_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_ec_rst_2.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_ec_rst_2.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_ec_rst_2.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_ec_rst_2.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_gsc_rst_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_gsc_rst_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_gsc_rst_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_gsc_rst_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_interrupt_2.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_interrupt_2.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_interrupt_2.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_interrupt_2.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_bat_disable_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_bat_disable_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_bat_disable_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_bat_disable_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_ec_rst_3.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_ec_rst_3.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_ec_rst_3.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_ec_rst_3.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_gsc_rst_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_gsc_rst_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_gsc_rst_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_gsc_rst_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_interrupt_3.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_interrupt_3.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_interrupt_3.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_interrupt_3.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_ac_present_sel_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_ac_present_sel_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_ac_present_sel_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_ac_present_sel_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key0_in_sel_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key0_in_sel_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key0_in_sel_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key0_in_sel_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key1_in_sel_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key1_in_sel_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key1_in_sel_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key1_in_sel_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key2_in_sel_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key2_in_sel_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key2_in_sel_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key2_in_sel_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_pwrb_in_sel_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_pwrb_in_sel_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_pwrb_in_sel_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_pwrb_in_sel_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_ac_present_sel_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_ac_present_sel_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_ac_present_sel_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_ac_present_sel_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key0_in_sel_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key0_in_sel_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key0_in_sel_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key0_in_sel_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key1_in_sel_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key1_in_sel_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key1_in_sel_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key1_in_sel_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key2_in_sel_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key2_in_sel_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key2_in_sel_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key2_in_sel_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_pwrb_in_sel_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_pwrb_in_sel_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_pwrb_in_sel_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_pwrb_in_sel_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_ac_present_sel_2.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_ac_present_sel_2.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_ac_present_sel_2.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_ac_present_sel_2.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key0_in_sel_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key0_in_sel_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key0_in_sel_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key0_in_sel_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key1_in_sel_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key1_in_sel_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key1_in_sel_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key1_in_sel_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key2_in_sel_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key2_in_sel_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key2_in_sel_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key2_in_sel_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_pwrb_in_sel_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_pwrb_in_sel_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_pwrb_in_sel_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_pwrb_in_sel_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_ac_present_sel_3.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_ac_present_sel_3.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_ac_present_sel_3.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_ac_present_sel_3.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key0_in_sel_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key0_in_sel_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key0_in_sel_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key0_in_sel_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key1_in_sel_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key1_in_sel_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key1_in_sel_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key1_in_sel_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key2_in_sel_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key2_in_sel_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key2_in_sel_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key2_in_sel_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_pwrb_in_sel_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_pwrb_in_sel_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_pwrb_in_sel_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_pwrb_in_sel_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo0_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo0_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo0_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo0_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo1_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo1_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo1_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo1_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo2_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo2_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo2_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo2_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo3_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo3_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo3_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo3_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_ec_rst_ctl.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_ec_rst_ctl.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_ec_rst_ctl.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_ec_rst_ctl.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_intr_enable.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_intr_enable.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_intr_enable.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_intr_enable.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_intr_state.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_intr_state.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_intr_state.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_intr_state.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_h2l.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_h2l.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_h2l.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_h2l.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_l2h.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_l2h.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_l2h.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_l2h.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_h2l.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_h2l.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_h2l.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_h2l.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_l2h.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_l2h.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_l2h.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_l2h.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_debounce_ctl.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_debounce_ctl.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_debounce_ctl.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_debounce_ctl.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_h2l.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_h2l.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_h2l.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_h2l.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_l2h.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_l2h.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_l2h.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_l2h.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_h2l.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_h2l.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_h2l.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_h2l.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_l2h.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_l2h.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_l2h.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_l2h.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_h2l.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_h2l.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_h2l.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_h2l.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_l2h.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_l2h.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_l2h.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_l2h.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_h2l.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_h2l.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_h2l.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_h2l.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_l2h.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_l2h.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_l2h.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_l2h.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_ac_present.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_ac_present.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_ac_present.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_ac_present.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_bat_disable.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_bat_disable.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_bat_disable.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_bat_disable.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_in.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_in.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_in.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_in.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_out.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_out.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_out.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_out.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_in.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_in.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_in.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_in.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_out.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_out.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_out.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_out.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_in.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_in.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_in.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_in.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_out.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_out.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_out.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_out.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_in.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_in.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_in.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_in.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_out.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_out.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_out.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_out.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_0.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_0.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_0.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_0.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_1.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_1.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_1.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_1.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ac_present.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ac_present.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ac_present.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ac_present.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ec_rst_l.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ec_rst_l.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ec_rst_l.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ec_rst_l.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key0_in.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key0_in.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key0_in.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key0_in.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key1_in.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key1_in.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key1_in.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key1_in.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key2_in.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key2_in.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key2_in.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key2_in.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_pwrb_in.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_pwrb_in.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_pwrb_in.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_pwrb_in.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_bat_disable.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_bat_disable.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_bat_disable.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_bat_disable.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_ec_rst_l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_ec_rst_l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_ec_rst_l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_ec_rst_l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key0_out.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key0_out.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key0_out.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key0_out.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key1_out.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key1_out.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key1_out.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key1_out.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key2_out.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key2_out.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key2_out.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key2_out.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_pwrb_out.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_pwrb_out.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_pwrb_out.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_pwrb_out.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_bat_disable.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_bat_disable.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_bat_disable.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_bat_disable.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_ec_rst_l.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_ec_rst_l.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_ec_rst_l.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_ec_rst_l.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key0_out.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key0_out.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key0_out.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key0_out.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key1_out.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key1_out.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key1_out.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key1_out.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key2_out.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key2_out.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key2_out.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key2_out.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_pwrb_out.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_pwrb_out.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_pwrb_out.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_pwrb_out.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_regwen.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_regwen.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_regwen.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.intg_error_q == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.intg_error_q  &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_llpbk.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_llpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_llpbk.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_llpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_nco.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_nco.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_nco.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_nco.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_nf.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_nf.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_nf.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_nf.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_parity_en.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_parity_en.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_parity_en.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_parity_en.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_parity_odd.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_parity_odd.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_parity_odd.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_parity_odd.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_rx.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_rx.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_rx.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_rx.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_rxblvl.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_rxblvl.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_rxblvl.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_rxblvl.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_slpbk.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_slpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_slpbk.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_slpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_tx.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_tx.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_tx.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_tx.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_rxilvl.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_rxilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_rxilvl.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_rxilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_rxrst.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_rxrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_rxrst.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_rxrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_txilvl.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_txilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_txilvl.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_txilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_txrst.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_txrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_txrst.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_txrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_break_err.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_break_err.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_break_err.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_break_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_frame_err.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_frame_err.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_frame_err.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_frame_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_overflow.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_overflow.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_parity_err.q   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_parity_err.q    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_parity_err.qe  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_parity_err.qe   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_timeout.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_timeout.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_tx_empty.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_tx_empty.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_tx_empty.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_tx_empty.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_break_err.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_break_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_break_err.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_break_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_frame_err.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_frame_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_frame_err.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_frame_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_parity_err.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_parity_err.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_parity_err.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_parity_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_timeout.q   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_timeout.qe  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_watermark.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_tx_empty.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_tx_watermark.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_tx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_tx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_tx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ovrd_txen.q   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ovrd_txen.q    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ovrd_txen.qe  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ovrd_txen.qe   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ovrd_txval.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ovrd_txval.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ovrd_txval.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ovrd_txval.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_timeout_ctrl_en.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_timeout_ctrl_en.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_timeout_ctrl_en.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_timeout_ctrl_en.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_timeout_ctrl_val.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_timeout_ctrl_val.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_timeout_ctrl_val.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_timeout_ctrl_val.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_wdata.q   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_wdata.q    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_wdata.qe  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_wdata.qe   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.allzero_cnt_q   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.allzero_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.break_st_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.break_st_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_break_err.intr_o == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_break_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_frame_err.intr_o == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_frame_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_overflow.intr_o  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_overflow.intr_o   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_parity_err.intr_o    == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_parity_err.intr_o &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_tx_empty.intr_o == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_tx_empty.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_tx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_tx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.nco_sum_q   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.nco_sum_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_fifo_depth_prev_q    == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_fifo_depth_prev_q &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_sync_q1  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_sync_q1   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_sync_q2  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_sync_q2   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_timeout_count_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_timeout_count_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_val_q    == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_val_q &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.tx_out_q    == top_level_upec.top_earlgrey_2.u_uart0.uart_core.tx_out_q &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.tx_uart_idle_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.tx_uart_idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.tx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart0.uart_core.tx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.idle_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.rx_valid_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.rx_valid_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_tx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_tx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_tx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_tx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_tx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_tx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_tx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_tx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_tx.tx_q    == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_tx.tx_q &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_llpbk.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_llpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_llpbk.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_llpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_nco.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_nco.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_nco.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_nco.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_nf.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_nf.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_nf.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_nf.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_parity_en.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_parity_en.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_parity_en.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_parity_en.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_parity_odd.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_parity_odd.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_parity_odd.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_parity_odd.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_rx.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_rx.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_rx.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_rx.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_rxblvl.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_rxblvl.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_rxblvl.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_rxblvl.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_slpbk.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_slpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_slpbk.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_slpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_tx.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_tx.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_tx.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_tx.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_rxilvl.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_rxilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_rxilvl.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_rxilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_rxrst.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_rxrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_rxrst.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_rxrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_txilvl.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_txilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_txilvl.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_txilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_txrst.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_txrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_txrst.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_txrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_break_err.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_break_err.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_break_err.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_break_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_frame_err.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_frame_err.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_frame_err.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_frame_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_overflow.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_overflow.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_parity_err.q   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_parity_err.q    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_parity_err.qe  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_parity_err.qe   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_timeout.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_timeout.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_tx_empty.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_tx_empty.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_tx_empty.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_tx_empty.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_break_err.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_break_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_break_err.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_break_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_frame_err.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_frame_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_frame_err.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_frame_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_parity_err.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_parity_err.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_parity_err.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_parity_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_timeout.q   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_timeout.qe  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_watermark.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_tx_empty.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_tx_watermark.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_tx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_tx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_tx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ovrd_txen.q   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ovrd_txen.q    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ovrd_txen.qe  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ovrd_txen.qe   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ovrd_txval.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ovrd_txval.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ovrd_txval.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ovrd_txval.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_timeout_ctrl_en.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_timeout_ctrl_en.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_timeout_ctrl_en.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_timeout_ctrl_en.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_timeout_ctrl_val.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_timeout_ctrl_val.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_timeout_ctrl_val.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_timeout_ctrl_val.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_wdata.q   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_wdata.q    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_wdata.qe  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_wdata.qe   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.allzero_cnt_q   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.allzero_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.break_st_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.break_st_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_break_err.intr_o == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_break_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_frame_err.intr_o == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_frame_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_overflow.intr_o  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_overflow.intr_o   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_parity_err.intr_o    == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_parity_err.intr_o &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_tx_empty.intr_o == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_tx_empty.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_tx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_tx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.nco_sum_q   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.nco_sum_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_fifo_depth_prev_q    == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_fifo_depth_prev_q &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_sync_q1  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_sync_q1   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_sync_q2  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_sync_q2   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_timeout_count_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_timeout_count_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_val_q    == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_val_q &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.tx_out_q    == top_level_upec.top_earlgrey_2.u_uart1.uart_core.tx_out_q &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.tx_uart_idle_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.tx_uart_idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.tx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart1.uart_core.tx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.idle_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.rx_valid_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.rx_valid_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_tx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_tx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_tx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_tx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_tx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_tx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_tx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_tx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_tx.tx_q    == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_tx.tx_q &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_llpbk.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_llpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_llpbk.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_llpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_nco.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_nco.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_nco.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_nco.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_nf.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_nf.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_nf.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_nf.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_parity_en.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_parity_en.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_parity_en.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_parity_en.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_parity_odd.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_parity_odd.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_parity_odd.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_parity_odd.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_rx.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_rx.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_rx.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_rx.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_rxblvl.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_rxblvl.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_rxblvl.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_rxblvl.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_slpbk.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_slpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_slpbk.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_slpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_tx.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_tx.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_tx.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_tx.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_rxilvl.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_rxilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_rxilvl.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_rxilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_rxrst.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_rxrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_rxrst.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_rxrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_txilvl.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_txilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_txilvl.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_txilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_txrst.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_txrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_txrst.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_txrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_break_err.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_break_err.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_break_err.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_break_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_frame_err.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_frame_err.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_frame_err.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_frame_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_overflow.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_overflow.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_parity_err.q   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_parity_err.q    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_parity_err.qe  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_parity_err.qe   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_timeout.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_timeout.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_tx_empty.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_tx_empty.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_tx_empty.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_tx_empty.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_break_err.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_break_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_break_err.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_break_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_frame_err.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_frame_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_frame_err.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_frame_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_parity_err.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_parity_err.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_parity_err.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_parity_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_timeout.q   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_timeout.qe  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_watermark.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_tx_empty.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_tx_watermark.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_tx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_tx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_tx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ovrd_txen.q   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ovrd_txen.q    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ovrd_txen.qe  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ovrd_txen.qe   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ovrd_txval.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ovrd_txval.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ovrd_txval.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ovrd_txval.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_timeout_ctrl_en.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_timeout_ctrl_en.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_timeout_ctrl_en.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_timeout_ctrl_en.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_timeout_ctrl_val.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_timeout_ctrl_val.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_timeout_ctrl_val.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_timeout_ctrl_val.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_wdata.q   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_wdata.q    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_wdata.qe  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_wdata.qe   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.allzero_cnt_q   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.allzero_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.break_st_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.break_st_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_break_err.intr_o == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_break_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_frame_err.intr_o == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_frame_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_overflow.intr_o  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_overflow.intr_o   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_parity_err.intr_o    == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_parity_err.intr_o &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_tx_empty.intr_o == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_tx_empty.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_tx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_tx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.nco_sum_q   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.nco_sum_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_fifo_depth_prev_q    == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_fifo_depth_prev_q &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_sync_q1  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_sync_q1   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_sync_q2  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_sync_q2   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_timeout_count_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_timeout_count_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_val_q    == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_val_q &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.tx_out_q    == top_level_upec.top_earlgrey_2.u_uart2.uart_core.tx_out_q &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.tx_uart_idle_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.tx_uart_idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.tx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart2.uart_core.tx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.idle_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.rx_valid_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.rx_valid_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_tx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_tx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_tx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_tx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_tx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_tx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_tx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_tx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_tx.tx_q    == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_tx.tx_q &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_llpbk.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_llpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_llpbk.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_llpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_nco.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_nco.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_nco.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_nco.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_nf.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_nf.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_nf.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_nf.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_parity_en.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_parity_en.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_parity_en.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_parity_en.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_parity_odd.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_parity_odd.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_parity_odd.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_parity_odd.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_rx.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_rx.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_rx.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_rx.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_rxblvl.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_rxblvl.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_rxblvl.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_rxblvl.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_slpbk.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_slpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_slpbk.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_slpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_tx.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_tx.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_tx.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_tx.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_rxilvl.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_rxilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_rxilvl.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_rxilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_rxrst.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_rxrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_rxrst.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_rxrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_txilvl.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_txilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_txilvl.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_txilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_txrst.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_txrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_txrst.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_txrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_break_err.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_break_err.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_break_err.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_break_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_frame_err.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_frame_err.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_frame_err.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_frame_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_overflow.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_overflow.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_parity_err.q   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_parity_err.q    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_parity_err.qe  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_parity_err.qe   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_timeout.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_timeout.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_tx_empty.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_tx_empty.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_tx_empty.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_tx_empty.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_break_err.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_break_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_break_err.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_break_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_frame_err.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_frame_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_frame_err.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_frame_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_parity_err.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_parity_err.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_parity_err.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_parity_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_timeout.q   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_timeout.qe  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_watermark.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_tx_empty.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_tx_watermark.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_tx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_tx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_tx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ovrd_txen.q   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ovrd_txen.q    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ovrd_txen.qe  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ovrd_txen.qe   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ovrd_txval.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ovrd_txval.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ovrd_txval.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ovrd_txval.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_timeout_ctrl_en.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_timeout_ctrl_en.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_timeout_ctrl_en.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_timeout_ctrl_en.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_timeout_ctrl_val.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_timeout_ctrl_val.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_timeout_ctrl_val.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_timeout_ctrl_val.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_wdata.q   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_wdata.q    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_wdata.qe  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_wdata.qe   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.allzero_cnt_q   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.allzero_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.break_st_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.break_st_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_break_err.intr_o == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_break_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_frame_err.intr_o == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_frame_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_overflow.intr_o  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_overflow.intr_o   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_parity_err.intr_o    == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_parity_err.intr_o &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_tx_empty.intr_o == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_tx_empty.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_tx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_tx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.nco_sum_q   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.nco_sum_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_fifo_depth_prev_q    == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_fifo_depth_prev_q &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_sync_q1  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_sync_q1   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_sync_q2  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_sync_q2   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_timeout_count_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_timeout_count_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_val_q    == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_val_q &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.tx_out_q    == top_level_upec.top_earlgrey_2.u_uart3.uart_core.tx_out_q &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.tx_uart_idle_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.tx_uart_idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.tx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart3.uart_core.tx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.idle_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.rx_valid_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.rx_valid_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_tx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_tx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_tx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_tx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_tx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_tx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_tx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_tx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_tx.tx_q    == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_tx.tx_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.aon_tgl  == top_level_upec.top_earlgrey_2.u_usbdev.aon_tgl   &&
        top_level_upec.top_earlgrey_1.u_usbdev.cdc_sys_to_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.cdc_sys_to_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.cdc_sys_to_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.cdc_sys_to_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.cdc_usb_to_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.cdc_usb_to_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.cdc_usb_to_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.cdc_usb_to_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.event_link_reset_q   == top_level_upec.top_earlgrey_2.u_usbdev.event_link_reset_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.i_usbdev_iomux.cdc_io_to_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.i_usbdev_iomux.cdc_io_to_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.i_usbdev_iomux.cdc_io_to_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.i_usbdev_iomux.cdc_io_to_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.i_usbdev_iomux.cdc_io_to_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.i_usbdev_iomux.cdc_io_to_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.i_usbdev_iomux.cdc_io_to_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.i_usbdev_iomux.cdc_io_to_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_av_empty.intr_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_av_empty.intr_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_av_overflow.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_av_overflow.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_connected.intr_o    == top_level_upec.top_earlgrey_2.u_usbdev.intr_connected.intr_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_disconnected.intr_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_disconnected.intr_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_frame.intr_o    == top_level_upec.top_earlgrey_2.u_usbdev.intr_frame.intr_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_host_lost.intr_o    == top_level_upec.top_earlgrey_2.u_usbdev.intr_host_lost.intr_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_hw_pkt_received.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_hw_pkt_received.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_hw_pkt_sent.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_hw_pkt_sent.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_in_err.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_in_err.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_out_err.intr_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_out_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_reset.intr_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_reset.intr_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_resume.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_resume.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_suspend.intr_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_suspend.intr_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_bitstuff_err.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_bitstuff_err.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_crc_err.intr_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_crc_err.intr_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_full.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_full.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_pid_err.intr_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_pid_err.intr_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_av_empty.dst_level_q  == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_av_empty.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_av_empty.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_av_empty.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_av_empty.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_av_empty.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_av_empty.src_level    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_av_empty.src_level &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_frame.dst_level_q == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_frame.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_frame.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_frame.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_frame.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_frame.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_frame.src_level   == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_frame.src_level    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_bitstuff_err.dst_level_q   == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_bitstuff_err.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_bitstuff_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_bitstuff_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_bitstuff_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_bitstuff_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_bitstuff_err.src_level == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_bitstuff_err.src_level  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_crc_err.dst_level_q    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_crc_err.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_crc_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_crc_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_crc_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_crc_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_crc_err.src_level  == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_crc_err.src_level   &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_full.dst_level_q   == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_full.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_full.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_full.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_full.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_full.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_full.src_level == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_full.src_level  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_pid_err.dst_level_q    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_pid_err.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_pid_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_pid_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_pid_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_pid_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_pid_err.src_level  == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_pid_err.src_level   &&
        top_level_upec.top_earlgrey_1.u_usbdev.syncevent.d_sync_q   == top_level_upec.top_earlgrey_2.u_usbdev.syncevent.d_sync_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.syncevent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.syncevent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.syncevent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.syncevent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.tgl_sync_d1  == top_level_upec.top_earlgrey_2.u_usbdev.tgl_sync_d1   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.a_rvalid_sram_q  == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.a_rvalid_sram_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.b_rvalid_sram_q  == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.b_rvalid_sram_q   &&
      //  top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o   == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o    &&
     //   top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o   == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o    &&
     //   top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.mem == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.mem  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_avbuffer.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_avbuffer.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_avbuffer.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_avbuffer.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_buffer_0.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_buffer_0.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_buffer_0.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_buffer_0.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_pend_0.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_pend_0.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_pend_0.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_pend_0.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_rdy_0.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_rdy_0.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_rdy_0.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_rdy_0.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_size_0.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_size_0.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_size_0.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_size_0.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_buffer_10.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_buffer_10.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_buffer_10.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_buffer_10.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_pend_10.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_pend_10.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_pend_10.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_pend_10.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_rdy_10.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_rdy_10.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_rdy_10.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_rdy_10.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_size_10.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_size_10.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_size_10.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_size_10.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_buffer_11.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_buffer_11.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_buffer_11.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_buffer_11.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_pend_11.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_pend_11.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_pend_11.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_pend_11.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_rdy_11.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_rdy_11.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_rdy_11.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_rdy_11.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_size_11.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_size_11.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_size_11.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_size_11.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_buffer_1.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_buffer_1.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_buffer_1.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_buffer_1.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_pend_1.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_pend_1.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_pend_1.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_pend_1.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_rdy_1.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_rdy_1.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_rdy_1.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_rdy_1.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_size_1.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_size_1.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_size_1.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_size_1.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_buffer_2.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_buffer_2.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_buffer_2.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_buffer_2.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_pend_2.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_pend_2.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_pend_2.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_pend_2.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_rdy_2.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_rdy_2.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_rdy_2.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_rdy_2.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_size_2.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_size_2.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_size_2.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_size_2.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_buffer_3.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_buffer_3.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_buffer_3.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_buffer_3.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_pend_3.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_pend_3.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_pend_3.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_pend_3.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_rdy_3.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_rdy_3.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_rdy_3.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_rdy_3.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_size_3.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_size_3.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_size_3.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_size_3.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_buffer_4.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_buffer_4.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_buffer_4.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_buffer_4.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_pend_4.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_pend_4.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_pend_4.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_pend_4.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_rdy_4.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_rdy_4.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_rdy_4.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_rdy_4.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_size_4.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_size_4.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_size_4.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_size_4.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_buffer_5.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_buffer_5.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_buffer_5.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_buffer_5.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_pend_5.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_pend_5.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_pend_5.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_pend_5.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_rdy_5.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_rdy_5.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_rdy_5.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_rdy_5.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_size_5.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_size_5.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_size_5.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_size_5.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_buffer_6.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_buffer_6.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_buffer_6.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_buffer_6.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_pend_6.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_pend_6.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_pend_6.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_pend_6.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_rdy_6.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_rdy_6.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_rdy_6.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_rdy_6.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_size_6.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_size_6.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_size_6.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_size_6.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_buffer_7.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_buffer_7.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_buffer_7.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_buffer_7.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_pend_7.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_pend_7.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_pend_7.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_pend_7.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_rdy_7.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_rdy_7.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_rdy_7.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_rdy_7.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_size_7.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_size_7.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_size_7.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_size_7.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_buffer_8.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_buffer_8.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_buffer_8.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_buffer_8.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_pend_8.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_pend_8.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_pend_8.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_pend_8.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_rdy_8.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_rdy_8.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_rdy_8.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_rdy_8.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_size_8.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_size_8.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_size_8.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_size_8.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_buffer_9.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_buffer_9.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_buffer_9.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_buffer_9.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_pend_9.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_pend_9.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_pend_9.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_pend_9.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_rdy_9.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_rdy_9.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_rdy_9.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_rdy_9.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_size_9.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_size_9.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_size_9.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_size_9.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_0.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_0.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_0.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_0.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_1.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_1.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_1.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_1.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_10.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_10.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_10.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_10.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_11.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_11.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_11.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_11.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_2.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_2.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_2.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_2.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_3.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_3.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_3.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_3.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_4.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_4.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_4.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_4.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_5.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_5.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_5.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_5.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_6.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_6.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_6.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_6.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_7.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_7.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_7.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_7.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_8.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_8.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_8.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_8.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_9.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_9.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_9.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_9.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_0.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_0.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_0.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_0.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_1.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_1.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_1.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_1.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_10.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_10.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_10.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_10.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_11.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_11.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_11.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_11.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_2.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_2.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_2.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_2.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_3.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_3.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_3.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_3.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_4.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_4.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_4.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_4.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_5.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_5.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_5.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_5.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_6.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_6.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_6.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_6.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_7.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_7.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_7.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_7.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_8.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_8.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_8.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_8.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_9.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_9.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_9.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_9.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_av_empty.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_av_empty.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_av_empty.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_av_empty.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_av_overflow.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_av_overflow.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_av_overflow.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_av_overflow.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_connected.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_connected.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_connected.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_connected.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_disconnected.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_disconnected.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_disconnected.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_disconnected.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_frame.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_frame.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_frame.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_frame.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_host_lost.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_host_lost.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_host_lost.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_host_lost.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_in_err.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_in_err.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_in_err.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_in_err.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_out_err.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_out_err.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_out_err.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_out_err.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_reset.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_reset.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_reset.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_reset.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_resume.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_resume.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_resume.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_resume.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_suspend.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_suspend.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_suspend.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_suspend.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_pkt_received.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_pkt_received.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_pkt_received.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_pkt_received.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_pkt_sent.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_pkt_sent.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_pkt_sent.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_pkt_sent.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_bitstuff_err.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_bitstuff_err.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_bitstuff_err.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_bitstuff_err.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_crc_err.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_crc_err.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_crc_err.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_crc_err.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_full.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_full.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_full.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_full.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_pid_err.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_pid_err.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_pid_err.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_pid_err.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_av_empty.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_av_empty.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_av_empty.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_av_empty.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_av_overflow.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_av_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_av_overflow.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_av_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_connected.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_connected.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_connected.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_connected.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_disconnected.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_disconnected.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_disconnected.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_disconnected.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_frame.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_frame.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_frame.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_frame.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_host_lost.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_host_lost.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_host_lost.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_host_lost.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_in_err.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_in_err.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_in_err.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_in_err.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_out_err.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_out_err.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_out_err.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_out_err.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_reset.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_reset.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_reset.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_reset.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_resume.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_resume.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_resume.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_resume.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_suspend.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_suspend.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_suspend.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_suspend.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_pkt_received.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_pkt_received.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_pkt_received.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_pkt_received.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_pkt_sent.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_pkt_sent.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_pkt_sent.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_pkt_sent.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_bitstuff_err.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_bitstuff_err.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_bitstuff_err.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_bitstuff_err.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_crc_err.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_crc_err.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_crc_err.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_crc_err.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_full.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_full.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_full.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_full.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_pid_err.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_pid_err.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_pid_err.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_pid_err.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_0.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_0.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_0.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_0.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_1.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_1.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_1.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_1.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_10.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_10.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_10.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_10.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_11.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_11.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_11.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_11.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_2.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_2.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_2.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_2.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_3.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_3.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_3.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_3.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_4.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_4.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_4.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_4.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_5.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_5.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_5.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_5.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_6.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_6.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_6.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_6.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_7.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_7.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_7.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_7.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_8.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_8.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_8.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_8.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_9.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_9.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_9.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_9.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_eop_single_bit.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_eop_single_bit.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_eop_single_bit.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_eop_single_bit.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_override_pwr_sense_en.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_override_pwr_sense_en.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_override_pwr_sense_en.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_override_pwr_sense_en.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_override_pwr_sense_val.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_override_pwr_sense_val.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_override_pwr_sense_val.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_override_pwr_sense_val.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_pinflip.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_pinflip.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_pinflip.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_pinflip.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_rx_differential_mode.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_rx_differential_mode.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_rx_differential_mode.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_rx_differential_mode.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_tx_differential_mode.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_tx_differential_mode.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_tx_differential_mode.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_tx_differential_mode.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_tx_osc_test_mode.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_tx_osc_test_mode.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_tx_osc_test_mode.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_tx_osc_test_mode.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_usb_ref_disable.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_usb_ref_disable.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_usb_ref_disable.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_usb_ref_disable.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_d_o.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_d_o.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_d_o.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_d_o.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dn_o.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dn_o.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dn_o.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dn_o.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dn_pullup_en_o.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dn_pullup_en_o.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dn_pullup_en_o.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dn_pullup_en_o.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dp_o.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dp_o.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dp_o.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dp_o.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dp_pullup_en_o.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dp_pullup_en_o.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dp_pullup_en_o.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dp_pullup_en_o.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_en.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_en.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_en.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_en.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_oe_o.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_oe_o.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_oe_o.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_oe_o.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_se0_o.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_se0_o.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_se0_o.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_se0_o.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_suspend_o.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_suspend_o.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_suspend_o.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_suspend_o.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_tx_mode_se_o.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_tx_mode_se_o.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_tx_mode_se_o.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_tx_mode_se_o.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_0.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_0.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_0.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_0.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_1.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_1.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_1.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_1.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_10.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_10.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_10.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_10.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_11.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_11.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_11.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_11.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_2.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_2.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_2.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_2.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_3.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_3.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_3.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_3.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_4.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_4.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_4.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_4.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_5.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_5.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_5.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_5.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_6.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_6.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_6.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_6.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_7.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_7.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_7.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_7.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_8.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_8.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_8.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_8.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_9.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_9.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_9.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_9.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_0.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_0.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_0.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_0.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_1.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_1.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_1.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_1.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_10.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_10.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_10.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_10.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_11.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_11.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_11.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_11.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_2.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_2.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_2.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_2.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_3.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_3.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_3.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_3.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_4.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_4.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_4.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_4.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_5.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_5.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_5.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_5.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_6.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_6.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_6.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_6.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_7.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_7.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_7.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_7.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_8.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_8.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_8.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_8.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_9.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_9.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_9.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_9.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.dev_select_outstanding    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.dev_select_outstanding &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.err_resp.err_opcode   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.err_resp.err_opcode    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.err_resp.err_req_pending  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.err_resp.err_req_pending   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.err_resp.err_rsp_pending  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.err_resp.err_rsp_pending   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.err_resp.err_size == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.err_resp.err_size  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.err_resp.err_source   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.err_resp.err_source    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.num_req_outstanding   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.num_req_outstanding    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_0.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_0.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_0.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_0.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_1.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_1.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_1.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_1.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_10.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_10.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_10.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_10.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_11.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_11.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_11.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_11.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_2.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_2.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_2.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_2.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_3.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_3.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_3.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_3.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_4.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_4.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_4.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_4.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_5.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_5.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_5.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_5.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_6.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_6.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_6.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_6.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_7.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_7.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_7.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_7.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_8.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_8.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_8.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_8.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_9.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_9.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_9.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_9.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_usbctrl_device_address.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_usbctrl_device_address.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_usbctrl_device_address.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_usbctrl_device_address.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_usbctrl_enable.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_usbctrl_enable.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_usbctrl_enable.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_usbctrl_enable.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_config_wake_ack.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_config_wake_ack.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_config_wake_ack.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_config_wake_ack.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_config_wake_en.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_config_wake_en.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_config_wake_en.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_config_wake_en.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_debug.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_debug.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_debug.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_debug.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tgl_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.u_tgl_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tgl_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.u_tgl_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.intg_error_q == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.intg_error_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usb_out_of_rst_o == top_level_upec.top_earlgrey_2.u_usbdev.usb_out_of_rst_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usb_ref_val_q    == top_level_upec.top_earlgrey_2.u_usbdev.usb_ref_val_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.storage    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.storage &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_data_toggle_clear.dst_level_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_data_toggle_clear.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_data_toggle_clear.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_data_toggle_clear.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_data_toggle_clear.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_data_toggle_clear.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_data_toggle_clear.src_level   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_data_toggle_clear.src_level    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_devclr.dst_level_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_devclr.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_devclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_devclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_devclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_devclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_devclr.src_level  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_devclr.src_level   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.av_rready_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.av_rready_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.frame_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.frame_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.ns_cnt   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.ns_cnt    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.out_max_used_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.out_max_used_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.pkt_start_rd == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.pkt_start_rd  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.std_write_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.std_write_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.data_toggle_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.data_toggle_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.ep_impl_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.ep_impl_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_current_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_current_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_data_get_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_data_get_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_get_addr_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_get_addr_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_newpkt_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_newpkt_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_rollback_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_rollback_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_xfr_state    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_xfr_state &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.tx_data_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.tx_data_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.current_xfer_setup_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.current_xfer_setup_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.data_toggle_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.data_toggle_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.ep_impl_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.ep_impl_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.nak_out_transfer   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.nak_out_transfer    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_current_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_current_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_data_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_data_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_data_put_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_data_put_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_newpkt_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_newpkt_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_put_addr_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_put_addr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_setup_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_setup_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_xfr_state  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_xfr_state   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.addr_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.addr_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bit_phase_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bit_phase_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bitstuff_error_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bitstuff_error_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bitstuff_history_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bitstuff_history_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.crc16_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.crc16_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.crc5_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.crc5_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.diff_state_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.diff_state_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.endp_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.endp_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.frame_num_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.frame_num_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.full_pid_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.full_pid_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_history_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_history_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_state_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_state_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_state_qq == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_state_qq  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.packet_valid_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.packet_valid_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.rx_data_buffer_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.rx_data_buffer_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.token_payload_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.token_payload_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bit_count_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bit_count_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bit_history_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bit_history_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q2   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q2    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q3   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q3    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q4   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q4    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.byte_strobe_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.byte_strobe_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.crc16_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.crc16_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.data_payload_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.data_payload_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.data_shift_reg_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.data_shift_reg_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.dp_eop_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.dp_eop_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.oe_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.oe_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.oe_shift_reg_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.oe_shift_reg_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.out_state_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.out_state_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.pid_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.pid_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.se0_shift_reg_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.se0_shift_reg_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.state_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.state_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.tx_data_get_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.tx_data_get_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.usb_d_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.usb_d_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.usb_se0_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.usb_se0_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_pwr_sense.stored_value_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_pwr_sense.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_pwr_sense.stored_vector_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_pwr_sense.stored_vector_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_se0.stored_value_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_se0.stored_value_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_se0.stored_vector_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_se0.stored_vector_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.host_presence_timer   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.host_presence_timer    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_inac_state_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_inac_state_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_inac_timer_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_inac_timer_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_rst_state_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_rst_state_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_rst_timer_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_rst_timer_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_state_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_state_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.wdata    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.wdata &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_outrdyclr.dst_level_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_outrdyclr.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_outrdyclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_outrdyclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_outrdyclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_outrdyclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_outrdyclr.src_level   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_outrdyclr.src_level    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rdysync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rdysync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rdysync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rdysync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_resume.dst_level_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_resume.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_resume.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_resume.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_resume.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_resume.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_resume.src_level  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_resume.src_level   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.storage    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.storage &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_setsent.dst_level_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_setsent.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_setsent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_setsent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_setsent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_setsent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_setsent.src_level == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_setsent.src_level  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_ep_cfg.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_ep_cfg.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_ep_cfg.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_ep_cfg.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_in_err.dst_level_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_in_err.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_in_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_in_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_in_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_in_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_in_err.src_level == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_in_err.src_level  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_out_err.dst_level_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_out_err.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_out_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_out_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_out_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_out_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_out_err.src_level    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_out_err.src_level &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_phy_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_phy_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_phy_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_phy_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o
    );
endfunction

function automatic soc_state_equivalence_peri_devices();
    soc_state_equivalence_peri_devices = (
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn0_max_v == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn0_max_v  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn0_min_v == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn0_min_v  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn1_max_v == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn1_max_v  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn1_min_v == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_chn1_min_v  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_lp_sample_cnt  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_lp_sample_cnt   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_np_sample_cnt  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_np_sample_cnt   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_pwrup_time == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_pwrup_time  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_wakeup_time    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.cfg_wakeup_time &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[0].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[1].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[2].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[3].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[4].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[5].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[6].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn0_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_cond.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_max_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.gen_filter_sync[7].i_cfg_chn1_min_v.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.dst_level_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.src_level  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_done.src_level   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.adc_ctrl_match_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.adc_ctrl_match_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn0_val    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn0_val &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn0_val_we == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn0_val_we  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn1_val    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn1_val &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn1_val_we == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.chn1_val_we  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.fsm_state_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.fsm_state_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.lp_sample_cnt_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.lp_sample_cnt_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.np_sample_cnt_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.np_sample_cnt_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.pwrup_timer_cnt_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.pwrup_timer_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.trigger_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.trigger_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.wakeup_timer_cnt_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_fsm.wakeup_timer_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_adc_ctrl_intr_o.intr_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_adc_ctrl_intr_o.intr_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.dst_level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.src_level    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_sink_det.src_level &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.dst_level_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.src_level == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det.src_level  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.dst_level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.src_level    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_1a5_src_det_flip.src_level &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.dst_level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.src_level    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_3a0_sink_det.src_level &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.dst_level_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.src_level  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_discon.src_level   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.dst_level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.src_level    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_sink_det.src_level &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.dst_level_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.src_level == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det.src_level  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.dst_level_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.src_level    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_adc_ctrl_intr.i_cc_src_det_flip.src_level &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_adc_enable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_adc_enable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_adc_enable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_adc_enable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.storage == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.storage  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn0_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.storage == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.storage  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_chn1_val_intr.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_fsm_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_fsm_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_fsm_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_fsm_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en3.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en3.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en3.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en3.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en5.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en5.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en5.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en5.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en6.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en6.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en6.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en6.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en7.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en7.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en7.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_intr_en7.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_lp_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.storage    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.storage &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_np_sample_cnt.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_intr_en.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_intr_en.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_intr_en.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_intr_en.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_oneshot_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_gray_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_sync_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_rptr_sync_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_wptr_gray_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_wptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_wptr_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.fifo_wptr_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.storage   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.storage    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_pwrup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en3.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en3.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en3.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en3.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en5.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en5.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en5.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en5.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en6.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en6.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en6.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en6.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en7.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en7.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en7.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_en7.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_gray_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_sync_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_rptr_sync_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_wptr_gray_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_wptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_wptr_q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.fifo_wptr_q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.storage  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.storage   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_cfg_wakeup_time.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.dst_level_q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.src_level   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.i_adc_ctrl_core.i_oneshot_done.src_level    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_cond_0.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_cond_0.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_cond_0.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_cond_0.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_max_v_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_max_v_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_max_v_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_max_v_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_min_v_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_min_v_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_min_v_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_0_min_v_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_cond_1.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_cond_1.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_cond_1.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_cond_1.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_max_v_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_max_v_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_max_v_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_max_v_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_min_v_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_min_v_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_min_v_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_1_min_v_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_cond_2.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_cond_2.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_cond_2.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_cond_2.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_max_v_2.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_max_v_2.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_max_v_2.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_max_v_2.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_min_v_2.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_min_v_2.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_min_v_2.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_2_min_v_2.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_cond_3.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_cond_3.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_cond_3.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_cond_3.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_max_v_3.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_max_v_3.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_max_v_3.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_max_v_3.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_min_v_3.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_min_v_3.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_min_v_3.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_3_min_v_3.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_cond_4.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_cond_4.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_cond_4.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_cond_4.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_max_v_4.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_max_v_4.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_max_v_4.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_max_v_4.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_min_v_4.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_min_v_4.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_min_v_4.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_4_min_v_4.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_cond_5.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_cond_5.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_cond_5.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_cond_5.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_max_v_5.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_max_v_5.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_max_v_5.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_max_v_5.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_min_v_5.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_min_v_5.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_min_v_5.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_5_min_v_5.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_cond_6.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_cond_6.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_cond_6.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_cond_6.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_max_v_6.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_max_v_6.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_max_v_6.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_max_v_6.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_min_v_6.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_min_v_6.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_min_v_6.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_6_min_v_6.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_cond_7.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_cond_7.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_cond_7.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_cond_7.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_max_v_7.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_max_v_7.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_max_v_7.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_max_v_7.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_min_v_7.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_min_v_7.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_min_v_7.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn0_filter_ctl_7_min_v_7.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_cond_0.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_cond_0.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_cond_0.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_cond_0.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_max_v_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_max_v_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_max_v_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_max_v_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_min_v_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_min_v_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_min_v_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_0_min_v_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_cond_1.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_cond_1.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_cond_1.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_cond_1.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_max_v_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_max_v_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_max_v_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_max_v_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_min_v_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_min_v_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_min_v_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_1_min_v_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_cond_2.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_cond_2.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_cond_2.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_cond_2.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_max_v_2.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_max_v_2.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_max_v_2.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_max_v_2.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_min_v_2.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_min_v_2.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_min_v_2.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_2_min_v_2.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_cond_3.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_cond_3.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_cond_3.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_cond_3.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_max_v_3.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_max_v_3.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_max_v_3.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_max_v_3.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_min_v_3.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_min_v_3.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_min_v_3.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_3_min_v_3.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_cond_4.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_cond_4.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_cond_4.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_cond_4.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_max_v_4.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_max_v_4.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_max_v_4.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_max_v_4.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_min_v_4.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_min_v_4.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_min_v_4.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_4_min_v_4.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_cond_5.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_cond_5.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_cond_5.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_cond_5.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_max_v_5.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_max_v_5.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_max_v_5.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_max_v_5.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_min_v_5.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_min_v_5.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_min_v_5.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_5_min_v_5.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_cond_6.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_cond_6.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_cond_6.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_cond_6.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_max_v_6.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_max_v_6.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_max_v_6.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_max_v_6.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_min_v_6.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_min_v_6.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_min_v_6.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_6_min_v_6.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_cond_7.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_cond_7.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_cond_7.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_cond_7.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_max_v_7.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_max_v_7.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_max_v_7.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_max_v_7.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_min_v_7.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_min_v_7.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_min_v_7.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn1_filter_ctl_7_min_v_7.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_ext_0.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_ext_0.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_ext_0.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_ext_0.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_0.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_0.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_0.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_0.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_ext_0.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_ext_0.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_ext_0.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_0_adc_chn_value_intr_ext_0.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_ext_1.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_ext_1.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_ext_1.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_ext_1.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_1.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_1.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_1.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_1.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_ext_1.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_ext_1.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_ext_1.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_chn_val_1_adc_chn_value_intr_ext_1.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_adc_enable.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_adc_enable.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_adc_enable.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_adc_enable.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_oneshot_mode.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_oneshot_mode.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_oneshot_mode.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_en_ctl_oneshot_mode.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_fsm_rst.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_fsm_rst.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_fsm_rst.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_fsm_rst.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter0_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter0_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter0_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter0_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter1_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter1_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter1_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter1_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter2_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter2_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter2_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter2_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter3_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter3_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter3_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter3_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter4_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter4_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter4_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter4_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter5_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter5_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter5_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter5_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter6_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter6_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter6_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter6_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter7_en.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter7_en.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter7_en.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_chn0_1_filter7_en.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_oneshot_intr_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_oneshot_intr_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_oneshot_intr_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_ctl_oneshot_intr_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_sink_det.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_sink_det.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_sink_det.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_sink_det.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det_flip.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det_flip.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det_flip.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_1a5_src_det_flip.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_3a0_sink_det.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_3a0_sink_det.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_3a0_sink_det.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_3a0_sink_det.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_discon.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_discon.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_discon.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_discon.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_sink_det.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_sink_det.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_sink_det.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_sink_det.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det_flip.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det_flip.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det_flip.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_cc_src_det_flip.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_oneshot.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_oneshot.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_intr_status_oneshot.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_intr_status_oneshot.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_lp_sample_ctl.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_lp_sample_ctl.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_lp_sample_ctl.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_lp_sample_ctl.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_lp_mode.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_lp_mode.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_lp_mode.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_lp_mode.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_pwrup_time.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_pwrup_time.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_pwrup_time.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_pwrup_time.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_wakeup_time.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_wakeup_time.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_wakeup_time.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_pd_ctl_wakeup_time.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_sample_ctl.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_sample_ctl.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_sample_ctl.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_sample_ctl.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter0_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter0_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter0_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter0_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter1_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter1_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter1_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter1_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter2_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter2_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter2_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter2_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter3_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter3_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter3_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter3_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter4_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter4_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter4_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter4_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter5_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter5_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter5_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter5_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter6_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter6_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter6_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter6_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter7_en.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter7_en.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter7_en.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_ctl_chn0_1_filter7_en.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_sink_det.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_sink_det.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_sink_det.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_sink_det.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det_flip.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det_flip.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det_flip.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_1a5_src_det_flip.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_3a0_sink_det.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_3a0_sink_det.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_3a0_sink_det.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_3a0_sink_det.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_discon.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_discon.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_discon.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_discon.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_sink_det.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_sink_det.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_sink_det.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_sink_det.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det.q == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det.q  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det.qe    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det.qe &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det_flip.q    == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det_flip.q &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det_flip.qe   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_adc_wakeup_status_cc_src_det_flip.qe    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_intr_enable.q  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_intr_enable.q   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_intr_enable.qe == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_intr_enable.qe  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_intr_state.q   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_intr_state.q    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_intr_state.qe  == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_intr_state.qe   &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_adc_ctrl_aon.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_adc_ctrl_aon.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[0].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[0].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[10].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[10].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[11].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[11].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[12].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[12].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[13].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[13].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[14].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[14].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[15].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[15].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[16].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[16].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[17].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[17].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[18].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[18].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[19].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[19].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[1].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[1].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[20].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[20].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[21].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[21].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[22].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[22].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[23].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[23].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[24].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[24].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[25].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[25].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[26].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[26].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[27].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[27].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[28].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[28].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[29].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[29].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[2].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[2].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[30].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[30].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[31].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[31].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[32].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[32].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[33].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[33].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[34].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[34].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[35].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[35].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[36].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[36].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[37].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[37].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[38].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[38].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[39].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[39].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[3].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[3].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[40].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[40].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[41].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[41].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[42].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[42].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[43].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[43].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[44].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[44].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[45].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[45].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[46].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[46].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[47].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[47].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[48].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[48].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[49].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[49].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[4].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[4].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[50].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[50].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.ping_pending_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.ping_pending_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.diff_nq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.diff_nq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.diff_pq  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.state_q  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.gen_async.state_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.level_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_decode_alert.level_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_prim_generic_flop_ack.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_prim_generic_flop_ack.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[51].u_alert_receiver.u_prim_generic_flop_ping.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[51].u_alert_receiver.u_prim_generic_flop_ping.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[5].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[5].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[6].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[6].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[7].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[7].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[8].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[8].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.ping_pending_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.ping_pending_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.ping_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.ping_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.state_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.state_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.u_decode_alert.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.u_decode_alert.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.u_decode_alert.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.u_prim_generic_flop_ack.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.u_prim_generic_flop_ack.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_alerts[9].u_alert_receiver.u_prim_generic_flop_ping.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_alerts[9].u_alert_receiver.u_prim_generic_flop_ping.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[0].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[0].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[0].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[0].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[0].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[0].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[0].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[0].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[0].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[0].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[1].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[1].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[1].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[1].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[1].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[1].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[1].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[1].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[1].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[1].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[2].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[2].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[2].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[2].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[2].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[2].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[2].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[2].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[2].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[2].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[3].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[3].u_accu.gen_double_accu[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[3].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[3].u_accu.gen_double_accu[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[3].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[3].u_esc_timer.gen_double_cnt[0].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[3].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[3].u_esc_timer.gen_double_cnt[1].u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_classes[3].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_classes[3].u_esc_timer.u_state_regs.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.esc_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.esc_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.esc_req_q1    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.esc_req_q1 &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.u_decode_resp.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.u_decode_resp.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[0].u_esc_sender.u_decode_resp.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[0].u_esc_sender.u_decode_resp.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.esc_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.esc_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.esc_req_q1    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.esc_req_q1 &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.u_decode_resp.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.u_decode_resp.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[1].u_esc_sender.u_decode_resp.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[1].u_esc_sender.u_decode_resp.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.esc_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.esc_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.esc_req_q1    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.esc_req_q1 &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.u_decode_resp.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.u_decode_resp.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[2].u_esc_sender.u_decode_resp.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[2].u_esc_sender.u_decode_resp.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.esc_req_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.esc_req_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.esc_req_q1    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.esc_req_q1 &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.ping_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.ping_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.state_q   == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.u_decode_resp.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.u_decode_resp.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_alert_handler.gen_esc_sev[3].u_esc_sender.u_decode_resp.level_q == top_level_upec.top_earlgrey_2.u_alert_handler.gen_esc_sev[3].u_esc_sender.u_decode_resp.level_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.fips_q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.fips_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_packer_fifo.clr_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_packer_fifo.clr_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_packer_fifo.data_q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_packer_fifo.data_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_packer_fifo.depth_q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_packer_fifo.depth_q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_packer_fifo.gen_unpack_mode.ptr_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_packer_fifo.gen_unpack_mode.ptr_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs   == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs   == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_cnt[0].u_prim_flop_en.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_cnt[0].u_prim_flop_en.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_cnt[1].u_prim_flop_en.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_cnt[1].u_prim_flop_en.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.cnt_q == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.perturbed_q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.perturbed_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.lfsr_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[0].u_prim_lfsr.lfsr_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.cnt_q == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.perturbed_q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.perturbed_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.lfsr_q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.gen_double_lfsr[1].u_prim_lfsr.lfsr_q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_ping_timer.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_alert_handler.u_ping_timer.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.i_irq_classa.intr_o    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.i_irq_classa.intr_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.i_irq_classb.intr_o    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.i_irq_classb.intr_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.i_irq_classc.intr_o    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.i_irq_classc.intr_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.i_irq_classd.intr_o    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.i_irq_classd.intr_o &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_10.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_10.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_10.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_10.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_11.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_11.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_11.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_11.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_12.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_12.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_12.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_12.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_13.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_13.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_13.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_13.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_14.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_14.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_14.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_14.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_15.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_15.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_15.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_15.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_16.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_16.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_16.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_16.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_17.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_17.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_17.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_17.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_18.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_18.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_18.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_18.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_19.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_19.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_19.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_19.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_20.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_20.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_20.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_20.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_21.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_21.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_21.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_21.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_22.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_22.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_22.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_22.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_23.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_23.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_23.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_23.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_24.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_24.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_24.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_24.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_25.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_25.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_25.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_25.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_26.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_26.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_26.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_26.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_27.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_27.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_27.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_27.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_28.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_28.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_28.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_28.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_29.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_29.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_29.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_29.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_30.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_30.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_30.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_30.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_31.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_31.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_31.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_31.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_32.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_32.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_32.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_32.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_33.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_33.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_33.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_33.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_34.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_34.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_34.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_34.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_35.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_35.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_35.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_35.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_36.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_36.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_36.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_36.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_37.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_37.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_37.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_37.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_38.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_38.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_38.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_38.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_39.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_39.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_39.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_39.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_4.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_4.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_4.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_4.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_40.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_40.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_40.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_40.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_41.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_41.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_41.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_41.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_42.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_42.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_42.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_42.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_43.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_43.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_43.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_43.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_44.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_44.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_44.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_44.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_45.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_45.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_45.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_45.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_46.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_46.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_46.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_46.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_47.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_47.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_47.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_47.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_48.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_48.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_48.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_48.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_49.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_49.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_49.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_49.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_5.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_5.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_5.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_5.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_50.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_50.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_50.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_50.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_51.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_51.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_51.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_51.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_6.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_6.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_6.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_6.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_7.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_7.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_7.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_7.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_8.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_8.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_8.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_8.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_9.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_9.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_9.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_cause_9.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_10.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_10.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_10.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_10.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_11.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_11.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_11.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_11.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_12.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_12.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_12.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_12.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_13.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_13.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_13.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_13.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_14.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_14.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_14.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_14.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_15.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_15.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_15.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_15.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_16.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_16.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_16.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_16.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_17.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_17.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_17.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_17.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_18.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_18.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_18.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_18.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_19.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_19.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_19.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_19.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_20.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_20.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_20.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_20.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_21.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_21.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_21.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_21.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_22.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_22.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_22.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_22.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_23.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_23.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_23.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_23.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_24.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_24.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_24.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_24.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_25.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_25.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_25.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_25.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_26.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_26.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_26.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_26.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_27.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_27.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_27.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_27.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_28.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_28.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_28.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_28.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_29.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_29.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_29.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_29.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_30.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_30.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_30.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_30.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_31.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_31.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_31.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_31.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_32.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_32.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_32.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_32.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_33.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_33.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_33.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_33.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_34.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_34.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_34.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_34.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_35.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_35.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_35.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_35.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_36.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_36.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_36.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_36.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_37.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_37.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_37.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_37.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_38.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_38.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_38.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_38.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_39.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_39.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_39.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_39.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_4.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_4.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_4.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_4.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_40.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_40.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_40.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_40.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_41.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_41.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_41.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_41.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_42.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_42.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_42.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_42.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_43.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_43.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_43.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_43.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_44.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_44.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_44.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_44.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_45.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_45.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_45.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_45.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_46.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_46.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_46.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_46.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_47.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_47.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_47.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_47.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_48.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_48.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_48.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_48.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_49.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_49.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_49.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_49.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_5.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_5.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_5.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_5.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_50.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_50.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_50.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_50.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_51.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_51.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_51.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_51.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_6.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_6.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_6.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_6.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_7.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_7.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_7.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_7.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_8.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_8.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_8.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_8.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_9.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_9.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_9.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_class_9.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_10.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_10.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_10.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_10.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_11.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_11.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_11.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_11.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_12.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_12.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_12.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_12.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_13.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_13.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_13.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_13.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_14.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_14.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_14.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_14.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_15.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_15.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_15.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_15.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_16.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_16.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_16.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_16.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_17.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_17.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_17.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_17.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_18.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_18.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_18.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_18.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_19.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_19.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_19.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_19.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_20.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_20.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_20.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_20.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_21.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_21.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_21.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_21.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_22.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_22.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_22.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_22.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_23.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_23.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_23.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_23.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_24.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_24.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_24.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_24.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_25.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_25.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_25.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_25.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_26.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_26.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_26.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_26.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_27.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_27.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_27.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_27.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_28.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_28.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_28.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_28.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_29.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_29.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_29.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_29.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_30.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_30.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_30.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_30.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_31.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_31.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_31.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_31.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_32.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_32.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_32.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_32.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_33.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_33.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_33.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_33.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_34.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_34.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_34.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_34.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_35.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_35.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_35.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_35.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_36.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_36.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_36.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_36.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_37.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_37.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_37.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_37.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_38.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_38.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_38.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_38.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_39.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_39.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_39.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_39.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_4.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_4.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_4.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_4.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_40.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_40.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_40.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_40.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_41.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_41.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_41.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_41.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_42.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_42.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_42.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_42.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_43.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_43.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_43.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_43.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_44.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_44.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_44.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_44.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_45.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_45.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_45.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_45.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_46.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_46.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_46.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_46.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_47.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_47.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_47.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_47.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_48.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_48.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_48.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_48.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_49.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_49.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_49.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_49.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_5.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_5.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_5.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_5.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_50.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_50.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_50.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_50.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_51.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_51.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_51.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_51.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_6.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_6.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_6.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_6.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_7.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_7.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_7.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_7.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_8.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_8.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_8.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_8.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_9.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_9.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_9.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_en_9.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_10.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_10.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_10.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_10.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_11.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_11.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_11.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_11.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_12.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_12.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_12.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_12.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_13.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_13.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_13.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_13.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_14.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_14.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_14.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_14.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_15.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_15.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_15.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_15.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_16.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_16.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_16.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_16.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_17.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_17.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_17.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_17.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_18.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_18.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_18.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_18.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_19.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_19.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_19.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_19.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_20.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_20.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_20.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_20.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_21.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_21.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_21.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_21.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_22.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_22.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_22.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_22.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_23.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_23.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_23.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_23.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_24.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_24.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_24.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_24.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_25.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_25.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_25.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_25.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_26.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_26.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_26.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_26.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_27.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_27.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_27.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_27.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_28.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_28.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_28.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_28.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_29.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_29.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_29.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_29.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_30.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_30.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_30.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_30.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_31.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_31.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_31.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_31.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_32.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_32.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_32.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_32.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_33.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_33.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_33.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_33.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_34.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_34.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_34.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_34.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_35.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_35.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_35.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_35.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_36.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_36.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_36.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_36.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_37.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_37.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_37.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_37.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_38.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_38.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_38.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_38.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_39.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_39.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_39.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_39.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_4.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_4.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_4.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_4.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_40.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_40.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_40.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_40.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_41.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_41.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_41.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_41.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_42.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_42.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_42.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_42.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_43.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_43.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_43.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_43.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_44.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_44.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_44.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_44.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_45.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_45.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_45.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_45.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_46.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_46.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_46.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_46.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_47.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_47.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_47.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_47.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_48.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_48.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_48.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_48.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_49.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_49.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_49.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_49.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_5.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_5.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_5.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_5.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_50.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_50.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_50.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_50.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_51.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_51.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_51.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_51.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_6.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_6.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_6.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_6.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_7.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_7.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_7.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_7.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_8.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_8.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_8.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_8.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_9.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_9.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_9.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_alert_regwen_9.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_accum_thresh.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_accum_thresh.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_accum_thresh.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_accum_thresh.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_clr_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_en_e3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_lock.q == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_lock.q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_lock.qe    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_lock.qe &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_ctrl_map_e3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase0_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase0_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase0_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase0_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase1_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase1_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase1_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase1_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase2_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase2_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase2_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase2_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase3_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase3_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase3_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_phase3_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_timeout_cyc.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_timeout_cyc.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classa_timeout_cyc.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classa_timeout_cyc.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_accum_thresh.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_accum_thresh.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_accum_thresh.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_accum_thresh.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_clr_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_en_e3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_lock.q == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_lock.q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_lock.qe    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_lock.qe &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_ctrl_map_e3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase0_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase0_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase0_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase0_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase1_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase1_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase1_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase1_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase2_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase2_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase2_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase2_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase3_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase3_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase3_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_phase3_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_timeout_cyc.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_timeout_cyc.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classb_timeout_cyc.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classb_timeout_cyc.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_accum_thresh.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_accum_thresh.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_accum_thresh.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_accum_thresh.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_clr_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_en_e3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_lock.q == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_lock.q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_lock.qe    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_lock.qe &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_ctrl_map_e3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase0_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase0_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase0_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase0_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase1_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase1_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase1_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase1_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase2_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase2_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase2_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase2_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase3_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase3_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase3_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_phase3_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_timeout_cyc.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_timeout_cyc.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classc_timeout_cyc.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classc_timeout_cyc.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_accum_thresh.q  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_accum_thresh.q   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_accum_thresh.qe == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_accum_thresh.qe  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_clr_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_en_e3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_lock.q == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_lock.q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_lock.qe    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_lock.qe &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_ctrl_map_e3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase0_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase0_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase0_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase0_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase1_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase1_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase1_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase1_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase2_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase2_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase2_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase2_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase3_cyc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase3_cyc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase3_cyc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_phase3_cyc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_timeout_cyc.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_timeout_cyc.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_classd_timeout_cyc.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_classd_timeout_cyc.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classa.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classa.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classa.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classa.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classb.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classb.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classb.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classb.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classc.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classc.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classc.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classc.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classd.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classd.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classd.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_enable_classd.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classa.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classa.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classa.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classa.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classb.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classb.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classb.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classb.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classc.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classc.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classc.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classc.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classd.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classd.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classd.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_intr_state_classd.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_4.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_4.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_4.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_cause_4.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_0.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_0.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_0.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_0.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_1.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_1.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_1.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_1.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_2.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_2.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_2.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_2.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_3.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_3.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_3.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_3.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_4.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_4.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_4.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_class_4.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_4.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_4.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_4.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_en_4.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_0.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_0.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_0.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_0.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_1.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_1.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_1.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_1.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_2.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_2.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_2.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_2.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_3.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_3.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_3.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_3.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_4.q   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_4.q    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_4.qe  == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_loc_alert_regwen_4.qe   &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timeout_cyc.q == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timeout_cyc.q  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timeout_cyc.qe    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timeout_cyc.qe &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_en.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_en.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_en.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_en.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_regwen.q    == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_regwen.q &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_regwen.qe   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_ping_timer_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_alert_handler.u_reg_wrap.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.aon_rst_req_q == top_level_upec.top_earlgrey_2.u_aon_timer_aon.aon_rst_req_q  &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.aon_wkup_req_q    == top_level_upec.top_earlgrey_2.u_aon_timer_aon.aon_wkup_req_q &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.prescale_count_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.prescale_count_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wdog_bark_thold_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wdog_bark_thold_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wdog_bite_thold_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wdog_bite_thold_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wdog_count_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wdog_count_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wdog_enable_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wdog_enable_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wdog_pause_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wdog_pause_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wkup_count_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wkup_count_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wkup_enable_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wkup_enable_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wkup_prescaler_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wkup_prescaler_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_core.wkup_thold_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_core.wkup_thold_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_intr_hw.intr_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_intr_hw.intr_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_intr_state_wdog_timer_expired.q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_intr_state_wdog_timer_expired.q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_intr_state_wdog_timer_expired.qe  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_intr_state_wdog_timer_expired.qe   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_intr_state_wkup_timer_expired.q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_intr_state_wkup_timer_expired.q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_intr_state_wkup_timer_expired.qe  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_intr_state_wkup_timer_expired.qe   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_wdog_regwen.q == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_wdog_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_reg.u_wdog_regwen.qe    == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_reg.u_wdog_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_sleep_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_sleep_mode.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_sleep_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_sleep_mode.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_wdog_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_wdog_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_wdog_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_wdog_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_wkup_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_wkup_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_sync_wkup_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_sync_wkup_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_gray_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_sync_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_rptr_sync_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_wptr_gray_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_wptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_wptr_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.fifo_wptr_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.storage   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.storage    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_gray_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_sync_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_rptr_sync_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_wptr_gray_q  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_wptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_wptr_q   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.fifo_wptr_q    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.storage   == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.storage    &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_aon_timer_aon.u_tlul_fifo.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.clk_status   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.clk_status    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.dis_status_q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.dis_status_q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.en_status_q  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.en_status_q   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div2_peri_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div2_peri_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div2_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div2_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div2_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div2_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div4_peri_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div4_peri_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div4_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div4_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_div4_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_div4_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_peri_cg.gen_generic.u_impl_generic.en_latch == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_peri_cg.gen_generic.u_impl_generic.en_latch  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_io_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_io_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_aes_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_aes_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_aes_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_aes_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_aes_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_aes_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_hmac_cg.gen_generic.u_impl_generic.en_latch   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_hmac_cg.gen_generic.u_impl_generic.en_latch    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_hmac_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_hmac_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_hmac_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_hmac_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_kmac_cg.gen_generic.u_impl_generic.en_latch   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_kmac_cg.gen_generic.u_impl_generic.en_latch    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_kmac_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_kmac_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_kmac_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_kmac_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_otbn_cg.gen_generic.u_impl_generic.en_latch   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_otbn_cg.gen_generic.u_impl_generic.en_latch    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_otbn_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_otbn_hint_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_main_otbn_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_main_otbn_hint_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_usb_peri_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_usb_peri_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_usb_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_usb_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clk_usb_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clk_usb_peri_sw_en_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clkmgr_byp.u_clk_byp_req.u_prim_flop.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clkmgr_byp.u_clk_byp_req.u_prim_flop.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clkmgr_byp.u_rcv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clkmgr_byp.u_rcv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clkmgr_byp.u_rcv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clkmgr_byp.u_rcv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_clkmgr_byp.u_send.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_clkmgr_byp.u_send.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_cg.i_cg.gen_generic.u_impl_generic.en_latch == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_cg.i_cg.gen_generic.u_impl_generic.en_latch  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div2_cg.i_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div2_cg.i_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div2_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div2_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div2_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div2_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div4_cg.i_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div4_cg.i_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div4_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div4_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_io_div4_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_io_div4_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_main_cg.i_cg.gen_generic.u_impl_generic.en_latch   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_main_cg.i_cg.gen_generic.u_impl_generic.en_latch    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_main_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_main_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_main_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_main_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_no_scan_io_div2_div.gen_div2.step_down_nq  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_no_scan_io_div2_div.gen_div2.step_down_nq   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_no_scan_io_div2_div.gen_div2.u_div2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_no_scan_io_div2_div.gen_div2.u_div2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_no_scan_io_div4_div.clk_int    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_no_scan_io_div4_div.clk_int &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_no_scan_io_div4_div.gen_div.cnt    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_no_scan_io_div4_div.gen_div.cnt &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_no_scan_io_div4_div.step_down_ack_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_no_scan_io_div4_div.step_down_ack_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div2_peri_en.q    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div2_peri_en.q &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div2_peri_en.qe   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div2_peri_en.qe    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div4_peri_en.q    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div4_peri_en.q &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div4_peri_en.qe   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_div4_peri_en.qe    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_peri_en.q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_peri_en.q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_peri_en.qe    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_io_peri_en.qe &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_usb_peri_en.q    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_usb_peri_en.q &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_enables_clk_usb_peri_en.qe   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_enables_clk_usb_peri_en.qe    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_aes_hint.q    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_aes_hint.q &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_aes_hint.qe   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_aes_hint.qe    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_hmac_hint.q   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_hmac_hint.q    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_hmac_hint.qe  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_hmac_hint.qe   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_kmac_hint.q   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_kmac_hint.q    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_kmac_hint.qe  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_kmac_hint.qe   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_otbn_hint.q   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_otbn_hint.q    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_otbn_hint.qe  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_clk_main_otbn_hint.qe   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_aes_val.q  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_aes_val.q   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_aes_val.qe == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_aes_val.qe  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_hmac_val.q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_hmac_val.q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_hmac_val.qe    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_hmac_val.qe &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_kmac_val.q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_kmac_val.q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_kmac_val.qe    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_kmac_val.qe &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_otbn_val.q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_otbn_val.q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_otbn_val.qe    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_clk_hints_status_clk_main_otbn_val.qe &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_extclk_sel.q == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_extclk_sel.q  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_extclk_sel.qe    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_extclk_sel.qe &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_extclk_sel_regwen.q  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_extclk_sel_regwen.q   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_extclk_sel_regwen.qe == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_extclk_sel_regwen.qe  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_jitter_enable.q  == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_jitter_enable.q   &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_jitter_enable.qe == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_jitter_enable.qe  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_roots_en_status_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_roots_en_status_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_roots_en_status_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_roots_en_status_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_roots_or_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_roots_or_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_roots_or_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_roots_or_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_usb_cg.i_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_usb_cg.i_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_usb_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_usb_cg.i_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_clkmgr_aon.u_usb_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_clkmgr_aon.u_usb_cg.i_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_gpio.cio_gpio_en_q  == top_level_upec.top_earlgrey_2.u_gpio.cio_gpio_en_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.cio_gpio_q == top_level_upec.top_earlgrey_2.u_gpio.cio_gpio_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.data_in_q  == top_level_upec.top_earlgrey_2.u_gpio.data_in_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_gpio.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[0].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[0].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[0].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[0].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[0].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[0].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[10].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[10].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[10].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[10].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[10].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[10].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[11].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[11].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[11].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[11].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[11].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[11].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[12].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[12].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[12].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[12].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[12].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[12].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[13].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[13].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[13].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[13].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[13].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[13].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[14].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[14].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[14].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[14].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[14].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[14].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[15].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[15].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[15].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[15].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[15].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[15].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[16].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[16].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[16].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[16].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[16].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[16].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[17].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[17].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[17].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[17].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[17].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[17].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[18].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[18].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[18].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[18].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[18].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[18].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[19].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[19].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[19].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[19].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[19].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[19].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[1].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[1].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[1].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[1].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[1].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[1].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[20].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[20].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[20].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[20].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[20].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[20].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[21].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[21].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[21].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[21].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[21].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[21].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[22].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[22].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[22].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[22].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[22].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[22].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[23].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[23].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[23].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[23].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[23].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[23].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[24].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[24].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[24].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[24].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[24].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[24].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[25].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[25].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[25].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[25].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[25].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[25].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[26].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[26].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[26].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[26].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[26].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[26].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[27].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[27].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[27].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[27].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[27].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[27].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[28].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[28].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[28].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[28].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[28].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[28].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[29].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[29].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[29].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[29].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[29].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[29].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[2].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[2].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[2].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[2].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[2].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[2].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[30].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[30].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[30].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[30].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[30].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[30].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[31].filter.diff_ctr_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[31].filter.diff_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[31].filter.filter_q == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[31].filter.filter_q  &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[31].filter.stored_value_q   == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[31].filter.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[3].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[3].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[3].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[3].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[3].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[3].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[4].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[4].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[4].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[4].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[4].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[4].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[5].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[5].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[5].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[5].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[5].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[5].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[6].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[6].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[6].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[6].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[6].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[6].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[7].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[7].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[7].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[7].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[7].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[7].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[8].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[8].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[8].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[8].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[8].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[8].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[9].filter.diff_ctr_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[9].filter.diff_ctr_q &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[9].filter.filter_q  == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[9].filter.filter_q   &&
        top_level_upec.top_earlgrey_1.u_gpio.gen_filter[9].filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_gpio.gen_filter[9].filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_gpio.intr_hw.intr_o == top_level_upec.top_earlgrey_2.u_gpio.intr_hw.intr_o  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_ctrl_en_input_filter.q == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_ctrl_en_input_filter.q  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_ctrl_en_input_filter.qe    == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_ctrl_en_input_filter.qe &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_data_in.q  == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_data_in.q   &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_data_in.qe == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_data_in.qe  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_falling.q == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_falling.q  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_falling.qe    == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_falling.qe &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_lvlhigh.q == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_lvlhigh.q  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_lvlhigh.qe    == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_lvlhigh.qe &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_lvllow.q  == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_lvllow.q   &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_lvllow.qe == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_lvllow.qe  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_rising.q  == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_rising.q   &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_ctrl_en_rising.qe == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_ctrl_en_rising.qe  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_enable.q  == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_enable.q   &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_enable.qe == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_enable.qe  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_state.q   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_state.q    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_intr_state.qe  == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_intr_state.qe   &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_gpio.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_gpio.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_i2c0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.fmt_watermark_q   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.fmt_watermark_q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_ack_stop.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_ack_stop.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_acq_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_acq_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_fmt_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_fmt_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_fmt_watermark.intr_o  == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_fmt_watermark.intr_o   &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_host_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_host_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_nak.intr_o    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_nak.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_rx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_rx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_rx_watermark.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_rx_watermark.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_scl_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_scl_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_sda_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_sda_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_sda_unstable.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_sda_unstable.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_stretch_timeout.intr_o    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_stretch_timeout.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_trans_complete.intr_o == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_trans_complete.intr_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_tx_empty.intr_o   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_tx_empty.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_tx_nonempty.intr_o    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_tx_nonempty.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.intr_hw_tx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.intr_hw_tx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.rx_watermark_q    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.rx_watermark_q &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.scl_rx_val    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.scl_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.sda_rx_val    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.sda_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.bit_idx == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.bit_idx  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.bit_index   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.bit_index    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.byte_index  == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.byte_index   &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.host_ack    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.host_ack &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.input_byte  == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.input_byte   &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.no_stop == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.no_stop  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.read_byte   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.read_byte    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.scl_high_cnt    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.scl_high_cnt &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.scl_i_q == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.scl_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.sda_i_q == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.sda_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.start_det   == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.start_det    &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.state_q == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.state_q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.stop_det    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.stop_det &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.stretch == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.stretch  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.stretch_stop_acq_clr    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.stretch_stop_acq_clr &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.stretch_stop_tx_clr == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.stretch_stop_tx_clr  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_fsm.tcount_q    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_fsm.tcount_q &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c0.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_enablehost.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_enablehost.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_enablehost.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_enablehost.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_enabletarget.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_enabletarget.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_enabletarget.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_enabletarget.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_llpbk.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_llpbk.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ctrl_llpbk.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ctrl_llpbk.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_fbyte.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_fbyte.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_fbyte.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_fbyte.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_nakok.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_nakok.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_nakok.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_nakok.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_rcont.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_rcont.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_rcont.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_rcont.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_read.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_read.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_read.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_read.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_start.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_start.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_start.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_start.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_stop.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_stop.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fdata_stop.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fdata_stop.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_acqrst.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_acqrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_acqrst.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_acqrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_fmtilvl.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_fmtilvl.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_fmtilvl.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_fmtilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_fmtrst.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_fmtrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_fmtrst.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_fmtrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_rxilvl.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_rxilvl.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_rxilvl.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_rxilvl.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_rxrst.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_rxrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_rxrst.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_rxrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_txrst.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_txrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_fifo_ctrl_txrst.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_fifo_ctrl_txrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_host_timeout_ctrl.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_host_timeout_ctrl.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_host_timeout_ctrl.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_host_timeout_ctrl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_ack_stop.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_ack_stop.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_ack_stop.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_ack_stop.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_acq_overflow.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_acq_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_acq_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_acq_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_fmt_overflow.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_fmt_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_fmt_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_fmt_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_fmt_watermark.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_fmt_watermark.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_fmt_watermark.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_fmt_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_host_timeout.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_host_timeout.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_host_timeout.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_host_timeout.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_nak.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_nak.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_nak.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_nak.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_rx_watermark.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_scl_interference.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_scl_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_scl_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_scl_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_sda_interference.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_sda_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_sda_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_sda_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_sda_unstable.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_sda_unstable.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_sda_unstable.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_sda_unstable.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_stretch_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_stretch_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_stretch_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_stretch_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_trans_complete.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_trans_complete.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_trans_complete.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_trans_complete.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_empty.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_nonempty.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_nonempty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_nonempty.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_nonempty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_enable_tx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_enable_tx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_ack_stop.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_ack_stop.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_ack_stop.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_ack_stop.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_acq_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_acq_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_acq_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_acq_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_fmt_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_fmt_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_fmt_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_fmt_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_fmt_watermark.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_fmt_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_fmt_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_fmt_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_host_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_host_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_host_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_host_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_nak.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_nak.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_nak.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_nak.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_rx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_rx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_rx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_rx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_rx_watermark.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_rx_watermark.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_rx_watermark.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_rx_watermark.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_scl_interference.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_scl_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_scl_interference.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_scl_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_sda_interference.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_sda_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_sda_interference.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_sda_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_sda_unstable.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_sda_unstable.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_sda_unstable.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_sda_unstable.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_stretch_timeout.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_stretch_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_stretch_timeout.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_stretch_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_trans_complete.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_trans_complete.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_trans_complete.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_trans_complete.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_empty.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_empty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_empty.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_empty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_nonempty.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_nonempty.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_nonempty.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_nonempty.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_intr_state_tx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_intr_state_tx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_sclval.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_sclval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_sclval.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_sclval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_sdaval.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_sdaval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_sdaval.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_sdaval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_txovrden.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_txovrden.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_ovrd_txovrden.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_ovrd_txovrden.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_en_addr_acq.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_en_addr_acq.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_en_addr_acq.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_en_addr_acq.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_en_addr_tx.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_en_addr_tx.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_en_addr_tx.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_en_addr_tx.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_stop_acq.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_stop_acq.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_stop_acq.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_stop_acq.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_stop_tx.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_stop_tx.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_stretch_ctrl_stop_tx.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_stretch_ctrl_stop_tx.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_address0.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_address0.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_address0.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_address0.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_address1.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_address1.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_address1.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_address1.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_mask0.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_mask0.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_mask0.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_mask0.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_mask1.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_mask1.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_target_id_mask1.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_target_id_mask1.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timeout_ctrl_en.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timeout_ctrl_en.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timeout_ctrl_en.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timeout_ctrl_en.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timeout_ctrl_val.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timeout_ctrl_val.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timeout_ctrl_val.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timeout_ctrl_val.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing0_thigh.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing0_thigh.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing0_thigh.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing0_thigh.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing0_tlow.q == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing0_tlow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing0_tlow.qe    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing0_tlow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing1_t_f.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing1_t_f.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing1_t_f.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing1_t_f.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing1_t_r.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing1_t_r.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing1_t_r.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing1_t_r.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing2_thd_sta.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing2_thd_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing2_thd_sta.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing2_thd_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing2_tsu_sta.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing2_tsu_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing2_tsu_sta.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing2_tsu_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing3_thd_dat.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing3_thd_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing3_thd_dat.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing3_thd_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing3_tsu_dat.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing3_tsu_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing3_tsu_dat.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing3_tsu_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing4_t_buf.q    == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing4_t_buf.q &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing4_t_buf.qe   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing4_t_buf.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing4_tsu_sto.q  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing4_tsu_sto.q   &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_timing4_tsu_sto.qe == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_timing4_tsu_sto.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_txdata.q   == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_txdata.q    &&
        top_level_upec.top_earlgrey_1.u_i2c0.u_reg.u_txdata.qe  == top_level_upec.top_earlgrey_2.u_i2c0.u_reg.u_txdata.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_i2c1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.fmt_watermark_q   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.fmt_watermark_q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_ack_stop.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_ack_stop.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_acq_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_acq_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_fmt_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_fmt_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_fmt_watermark.intr_o  == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_fmt_watermark.intr_o   &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_host_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_host_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_nak.intr_o    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_nak.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_rx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_rx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_rx_watermark.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_rx_watermark.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_scl_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_scl_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_sda_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_sda_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_sda_unstable.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_sda_unstable.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_stretch_timeout.intr_o    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_stretch_timeout.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_trans_complete.intr_o == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_trans_complete.intr_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_tx_empty.intr_o   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_tx_empty.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_tx_nonempty.intr_o    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_tx_nonempty.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.intr_hw_tx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.intr_hw_tx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.rx_watermark_q    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.rx_watermark_q &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.scl_rx_val    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.scl_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.sda_rx_val    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.sda_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.bit_idx == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.bit_idx  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.bit_index   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.bit_index    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.byte_index  == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.byte_index   &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.host_ack    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.host_ack &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.input_byte  == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.input_byte   &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.no_stop == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.no_stop  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.read_byte   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.read_byte    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.scl_high_cnt    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.scl_high_cnt &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.scl_i_q == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.scl_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.sda_i_q == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.sda_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.start_det   == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.start_det    &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.state_q == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.state_q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.stop_det    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.stop_det &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.stretch == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.stretch  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.stretch_stop_acq_clr    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.stretch_stop_acq_clr &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.stretch_stop_tx_clr == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.stretch_stop_tx_clr  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_fsm.tcount_q    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_fsm.tcount_q &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c1.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_enablehost.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_enablehost.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_enablehost.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_enablehost.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_enabletarget.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_enabletarget.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_enabletarget.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_enabletarget.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_llpbk.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_llpbk.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ctrl_llpbk.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ctrl_llpbk.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_fbyte.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_fbyte.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_fbyte.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_fbyte.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_nakok.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_nakok.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_nakok.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_nakok.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_rcont.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_rcont.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_rcont.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_rcont.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_read.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_read.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_read.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_read.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_start.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_start.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_start.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_start.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_stop.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_stop.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fdata_stop.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fdata_stop.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_acqrst.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_acqrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_acqrst.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_acqrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_fmtilvl.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_fmtilvl.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_fmtilvl.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_fmtilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_fmtrst.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_fmtrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_fmtrst.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_fmtrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_rxilvl.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_rxilvl.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_rxilvl.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_rxilvl.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_rxrst.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_rxrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_rxrst.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_rxrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_txrst.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_txrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_fifo_ctrl_txrst.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_fifo_ctrl_txrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_host_timeout_ctrl.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_host_timeout_ctrl.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_host_timeout_ctrl.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_host_timeout_ctrl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_ack_stop.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_ack_stop.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_ack_stop.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_ack_stop.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_acq_overflow.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_acq_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_acq_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_acq_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_fmt_overflow.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_fmt_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_fmt_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_fmt_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_fmt_watermark.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_fmt_watermark.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_fmt_watermark.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_fmt_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_host_timeout.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_host_timeout.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_host_timeout.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_host_timeout.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_nak.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_nak.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_nak.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_nak.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_rx_watermark.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_scl_interference.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_scl_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_scl_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_scl_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_sda_interference.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_sda_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_sda_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_sda_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_sda_unstable.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_sda_unstable.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_sda_unstable.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_sda_unstable.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_stretch_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_stretch_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_stretch_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_stretch_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_trans_complete.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_trans_complete.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_trans_complete.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_trans_complete.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_empty.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_nonempty.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_nonempty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_nonempty.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_nonempty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_enable_tx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_enable_tx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_ack_stop.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_ack_stop.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_ack_stop.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_ack_stop.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_acq_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_acq_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_acq_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_acq_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_fmt_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_fmt_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_fmt_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_fmt_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_fmt_watermark.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_fmt_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_fmt_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_fmt_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_host_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_host_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_host_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_host_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_nak.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_nak.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_nak.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_nak.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_rx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_rx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_rx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_rx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_rx_watermark.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_rx_watermark.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_rx_watermark.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_rx_watermark.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_scl_interference.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_scl_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_scl_interference.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_scl_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_sda_interference.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_sda_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_sda_interference.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_sda_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_sda_unstable.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_sda_unstable.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_sda_unstable.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_sda_unstable.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_stretch_timeout.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_stretch_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_stretch_timeout.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_stretch_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_trans_complete.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_trans_complete.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_trans_complete.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_trans_complete.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_empty.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_empty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_empty.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_empty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_nonempty.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_nonempty.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_nonempty.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_nonempty.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_intr_state_tx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_intr_state_tx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_sclval.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_sclval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_sclval.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_sclval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_sdaval.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_sdaval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_sdaval.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_sdaval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_txovrden.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_txovrden.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_ovrd_txovrden.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_ovrd_txovrden.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_en_addr_acq.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_en_addr_acq.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_en_addr_acq.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_en_addr_acq.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_en_addr_tx.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_en_addr_tx.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_en_addr_tx.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_en_addr_tx.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_stop_acq.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_stop_acq.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_stop_acq.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_stop_acq.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_stop_tx.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_stop_tx.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_stretch_ctrl_stop_tx.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_stretch_ctrl_stop_tx.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_address0.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_address0.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_address0.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_address0.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_address1.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_address1.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_address1.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_address1.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_mask0.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_mask0.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_mask0.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_mask0.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_mask1.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_mask1.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_target_id_mask1.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_target_id_mask1.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timeout_ctrl_en.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timeout_ctrl_en.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timeout_ctrl_en.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timeout_ctrl_en.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timeout_ctrl_val.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timeout_ctrl_val.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timeout_ctrl_val.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timeout_ctrl_val.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing0_thigh.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing0_thigh.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing0_thigh.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing0_thigh.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing0_tlow.q == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing0_tlow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing0_tlow.qe    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing0_tlow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing1_t_f.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing1_t_f.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing1_t_f.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing1_t_f.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing1_t_r.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing1_t_r.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing1_t_r.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing1_t_r.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing2_thd_sta.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing2_thd_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing2_thd_sta.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing2_thd_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing2_tsu_sta.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing2_tsu_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing2_tsu_sta.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing2_tsu_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing3_thd_dat.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing3_thd_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing3_thd_dat.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing3_thd_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing3_tsu_dat.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing3_tsu_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing3_tsu_dat.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing3_tsu_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing4_t_buf.q    == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing4_t_buf.q &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing4_t_buf.qe   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing4_t_buf.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing4_tsu_sto.q  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing4_tsu_sto.q   &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_timing4_tsu_sto.qe == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_timing4_tsu_sto.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_txdata.q   == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_txdata.q    &&
        top_level_upec.top_earlgrey_1.u_i2c1.u_reg.u_txdata.qe  == top_level_upec.top_earlgrey_2.u_i2c1.u_reg.u_txdata.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_i2c2.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.fmt_watermark_q   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.fmt_watermark_q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_ack_stop.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_ack_stop.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_acq_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_acq_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_fmt_overflow.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_fmt_overflow.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_fmt_watermark.intr_o  == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_fmt_watermark.intr_o   &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_host_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_host_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_nak.intr_o    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_nak.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_rx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_rx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_rx_watermark.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_rx_watermark.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_scl_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_scl_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_sda_interference.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_sda_interference.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_sda_unstable.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_sda_unstable.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_stretch_timeout.intr_o    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_stretch_timeout.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_trans_complete.intr_o == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_trans_complete.intr_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_tx_empty.intr_o   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_tx_empty.intr_o    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_tx_nonempty.intr_o    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_tx_nonempty.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.intr_hw_tx_overflow.intr_o    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.intr_hw_tx_overflow.intr_o &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.rx_watermark_q    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.rx_watermark_q &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.scl_rx_val    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.scl_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.sda_rx_val    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.sda_rx_val &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_acqfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fmtfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.bit_idx == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.bit_idx  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.bit_index   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.bit_index    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.byte_index  == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.byte_index   &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.host_ack    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.host_ack &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.input_byte  == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.input_byte   &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.no_stop == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.no_stop  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.read_byte   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.read_byte    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.scl_high_cnt    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.scl_high_cnt &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.scl_i_q == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.scl_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.sda_i_q == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.sda_i_q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.start_det   == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.start_det    &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.state_q == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.state_q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.stop_det    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.stop_det &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.stretch == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.stretch  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.stretch_stop_acq_clr    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.stretch_stop_acq_clr &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.stretch_stop_tx_clr == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.stretch_stop_tx_clr  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_fsm.tcount_q    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_fsm.tcount_q &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_rxfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_sync_scl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_sync_sda.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_i2c2.i2c_core.u_i2c_txfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_enablehost.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_enablehost.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_enablehost.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_enablehost.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_enabletarget.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_enabletarget.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_enabletarget.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_enabletarget.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_llpbk.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_llpbk.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ctrl_llpbk.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ctrl_llpbk.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_fbyte.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_fbyte.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_fbyte.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_fbyte.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_nakok.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_nakok.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_nakok.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_nakok.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_rcont.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_rcont.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_rcont.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_rcont.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_read.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_read.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_read.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_read.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_start.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_start.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_start.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_start.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_stop.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_stop.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fdata_stop.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fdata_stop.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_acqrst.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_acqrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_acqrst.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_acqrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_fmtilvl.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_fmtilvl.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_fmtilvl.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_fmtilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_fmtrst.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_fmtrst.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_fmtrst.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_fmtrst.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_rxilvl.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_rxilvl.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_rxilvl.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_rxilvl.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_rxrst.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_rxrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_rxrst.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_rxrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_txrst.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_txrst.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_fifo_ctrl_txrst.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_fifo_ctrl_txrst.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_host_timeout_ctrl.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_host_timeout_ctrl.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_host_timeout_ctrl.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_host_timeout_ctrl.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_ack_stop.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_ack_stop.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_ack_stop.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_ack_stop.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_acq_overflow.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_acq_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_acq_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_acq_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_fmt_overflow.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_fmt_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_fmt_overflow.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_fmt_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_fmt_watermark.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_fmt_watermark.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_fmt_watermark.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_fmt_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_host_timeout.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_host_timeout.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_host_timeout.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_host_timeout.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_nak.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_nak.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_nak.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_nak.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_rx_watermark.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_scl_interference.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_scl_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_scl_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_scl_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_sda_interference.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_sda_interference.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_sda_interference.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_sda_interference.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_sda_unstable.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_sda_unstable.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_sda_unstable.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_sda_unstable.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_stretch_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_stretch_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_stretch_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_stretch_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_trans_complete.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_trans_complete.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_trans_complete.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_trans_complete.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_empty.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_nonempty.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_nonempty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_nonempty.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_nonempty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_enable_tx_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_enable_tx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_ack_stop.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_ack_stop.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_ack_stop.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_ack_stop.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_acq_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_acq_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_acq_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_acq_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_fmt_overflow.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_fmt_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_fmt_overflow.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_fmt_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_fmt_watermark.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_fmt_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_fmt_watermark.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_fmt_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_host_timeout.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_host_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_host_timeout.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_host_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_nak.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_nak.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_nak.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_nak.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_rx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_rx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_rx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_rx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_rx_watermark.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_rx_watermark.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_rx_watermark.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_rx_watermark.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_scl_interference.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_scl_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_scl_interference.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_scl_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_sda_interference.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_sda_interference.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_sda_interference.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_sda_interference.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_sda_unstable.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_sda_unstable.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_sda_unstable.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_sda_unstable.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_stretch_timeout.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_stretch_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_stretch_timeout.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_stretch_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_trans_complete.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_trans_complete.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_trans_complete.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_trans_complete.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_empty.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_empty.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_empty.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_empty.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_nonempty.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_nonempty.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_nonempty.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_nonempty.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_overflow.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_intr_state_tx_overflow.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_intr_state_tx_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_sclval.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_sclval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_sclval.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_sclval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_sdaval.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_sdaval.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_sdaval.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_sdaval.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_txovrden.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_txovrden.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_ovrd_txovrden.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_ovrd_txovrden.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_en_addr_acq.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_en_addr_acq.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_en_addr_acq.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_en_addr_acq.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_en_addr_tx.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_en_addr_tx.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_en_addr_tx.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_en_addr_tx.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_stop_acq.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_stop_acq.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_stop_acq.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_stop_acq.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_stop_tx.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_stop_tx.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_stretch_ctrl_stop_tx.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_stretch_ctrl_stop_tx.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_address0.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_address0.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_address0.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_address0.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_address1.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_address1.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_address1.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_address1.qe   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_mask0.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_mask0.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_mask0.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_mask0.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_mask1.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_mask1.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_target_id_mask1.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_target_id_mask1.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timeout_ctrl_en.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timeout_ctrl_en.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timeout_ctrl_en.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timeout_ctrl_en.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timeout_ctrl_val.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timeout_ctrl_val.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timeout_ctrl_val.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timeout_ctrl_val.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing0_thigh.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing0_thigh.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing0_thigh.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing0_thigh.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing0_tlow.q == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing0_tlow.q  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing0_tlow.qe    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing0_tlow.qe &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing1_t_f.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing1_t_f.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing1_t_f.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing1_t_f.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing1_t_r.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing1_t_r.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing1_t_r.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing1_t_r.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing2_thd_sta.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing2_thd_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing2_thd_sta.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing2_thd_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing2_tsu_sta.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing2_tsu_sta.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing2_tsu_sta.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing2_tsu_sta.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing3_thd_dat.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing3_thd_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing3_thd_dat.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing3_thd_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing3_tsu_dat.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing3_tsu_dat.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing3_tsu_dat.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing3_tsu_dat.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing4_t_buf.q    == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing4_t_buf.q &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing4_t_buf.qe   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing4_t_buf.qe    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing4_tsu_sto.q  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing4_tsu_sto.q   &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_timing4_tsu_sto.qe == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_timing4_tsu_sto.qe  &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_txdata.q   == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_txdata.q    &&
        top_level_upec.top_earlgrey_1.u_i2c2.u_reg.u_txdata.qe  == top_level_upec.top_earlgrey_2.u_i2c2.u_reg.u_txdata.qe   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.fatal_bus_integ_error_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.fatal_bus_integ_error_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.fatal_prog_error_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.fatal_prog_error_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.fatal_state_error_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.fatal_state_error_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.flash_rma_error_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.flash_rma_error_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_set_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_set_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.ping_set_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.state_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.state_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_set_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_set_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_test_set_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_test_set_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.ping_set_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.ping_set_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.state_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.state_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.level_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.level_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.level_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.level_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_prim_generic_flop.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_prim_generic_flop.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.alert_set_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.alert_set_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.alert_test_set_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.alert_test_set_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.ping_set_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.ping_set_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.state_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.state_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ack.level_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ack.level_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ping.level_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_decode_ping.level_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_prim_generic_flop.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.gen_alert_tx[2].u_prim_alert_sender.u_prim_generic_flop.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_done_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_done_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.lc_idle_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.lc_idle_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.otp_part_error_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.otp_part_error_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.otp_test_ctrl_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.otp_test_ctrl_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.sw_claim_transition_if_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.sw_claim_transition_if_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.tap_claim_transition_if_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.tap_claim_transition_if_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.token_invalid_error_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.token_invalid_error_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.trans_cnt_oflw_error_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.trans_cnt_oflw_error_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.trans_invalid_error_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.trans_invalid_error_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.trans_success_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.trans_success_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.transition_target_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.transition_target_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.transition_token_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.transition_token_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.address_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.address_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.data_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.data_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.dr_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.dr_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.error_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.error_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_gray_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_sync_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_rptr_sync_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_wptr_gray_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_wptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_wptr_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.fifo_wptr_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.storage  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.storage   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_req.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.storage == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.storage  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_cdc.i_cdc_resp.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.bypass_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.bypass_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.dtmcs_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.dtmcs_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.idcode_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.idcode_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.jtag_ir_q == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.jtag_ir_q  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.jtag_ir_shift_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.jtag_ir_shift_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.tap_state_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.tap_state_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.td_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.td_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.tdo_oe_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.i_dmi_jtag_tap.tdo_oe_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_dmi_jtag.state_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_dmi_jtag.state_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.lc_state_valid_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.lc_state_valid_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_cnt_regs.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_cnt_regs.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_fsm_state_regs.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_fsm_state_regs.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_id_state_regs.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_id_state_regs.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_flo_keymgr_div.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_flo_keymgr_div.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_cpu_en.u_prim_flop.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_cpu_en.u_prim_flop.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_creator_seed_sw_rw_en.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_creator_seed_sw_rw_en.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_dft_en.u_prim_flop.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_dft_en.u_prim_flop.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_escalate_en.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_escalate_en.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_hw_debug_en.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_hw_debug_en.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_iso_part_sw_rd_en.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_iso_part_sw_rd_en.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_iso_part_sw_wr_en.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_iso_part_sw_wr_en.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_keymgr_en.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_keymgr_en.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_nvm_debug_en.u_prim_flop.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_nvm_debug_en.u_prim_flop.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_owner_seed_sw_rw_en.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_owner_seed_sw_rw_en.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_seed_hw_rd_en.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_seed_hw_rd_en.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_test_or_rma.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_lc_ctrl_signal_decode.u_prim_lc_sender_test_or_rma.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_check_byp_en.u_prim_flop.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_check_byp_en.u_prim_flop.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_clk_byp_req.u_prim_flop.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_clk_byp_req.u_prim_flop.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_flash_rma_req.u_prim_flop.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sender_flash_rma_req.u_prim_flop.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_clk_byp_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_clk_byp_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_clk_byp_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_clk_byp_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_flash_rma_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_flash_rma_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_flash_rma_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_prim_lc_sync_flash_rma_ack.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_fsm.u_state_regs.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_fsm.u_state_regs.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.hashed_token_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.hashed_token_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.token_hash_ack_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.token_hash_ack_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.token_hash_err_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.token_hash_err_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.gen_data_reg.data_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.gen_data_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.dst_ack_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.dst_ack_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.dst_fsm_cs  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.dst_fsm_cs   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.src_fsm_cs  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.src_fsm_cs   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.src_req_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_in.u_prim_sync_reqack.src_req_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.dst_ack_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.dst_ack_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.dst_fsm_cs == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.dst_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.src_fsm_cs == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.src_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.src_req_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_prim_sync_reqack_data_out.u_prim_sync_reqack.src_req_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_lc_ctrl_kmac_if.u_state_regs.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_lc_ctrl_kmac_if.u_state_regs.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver1.state_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver1.state_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver1.u_decode_esc.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver1.u_decode_esc.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver1.u_decode_esc.level_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver1.u_decode_esc.level_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver1.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver1.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver2.state_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver2.state_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver2.u_decode_esc.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver2.u_decode_esc.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver2.u_decode_esc.level_q   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver2.u_decode_esc.level_q    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_esc_receiver2.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_esc_receiver2.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_flop_2sync_init.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_flop_2sync_init.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_prim_flop_2sync_init.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_prim_flop_2sync_init.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.intg_err_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.intg_err_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_reg_tap.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_reg_tap.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_tap_tlul_host.g_multiple_reqs.source_q    == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_tap_tlul_host.g_multiple_reqs.source_q &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_tap_tlul_host.intg_err_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_tap_tlul_host.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_lc_ctrl.u_tap_tlul_host.outstanding_reqs_q  == top_level_upec.top_earlgrey_2.u_lc_ctrl.u_tap_tlul_host.outstanding_reqs_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.fatal_check_error_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.fatal_check_error_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.fatal_macro_error_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.fatal_macro_error_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_alert_tx[1].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.pending_tlul_error_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.pending_tlul_error_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.tlul_addr_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.tlul_addr_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[0].gen_unbuffered.u_part_unbuf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.pending_tlul_error_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.pending_tlul_error_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.tlul_addr_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.tlul_addr_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[1].gen_unbuffered.u_part_unbuf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.cnt_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.cnt_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.dout_gate_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.dout_gate_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[2].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.cnt_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.cnt_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.dout_gate_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.dout_gate_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[3].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.cnt_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.cnt_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.dout_gate_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.dout_gate_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[4].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.cnt_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.cnt_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.dout_gate_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.dout_gate_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.data_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[5].gen_buffered.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.cnt_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.cnt_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.dout_gate_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.dout_gate_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.error_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.error_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_otp_ctrl_ecc_reg.data_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_otp_ctrl_ecc_reg.data_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_otp_ctrl_ecc_reg.ecc_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.gen_partitions[6].gen_lifecycle.u_part_buf.u_state_regs.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.interrupt_triggers_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.interrupt_triggers_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.otp_idle_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.otp_idle_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.pwr_otp_rsp_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.pwr_otp_rsp_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.tlul_oob_err_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.tlul_oob_err_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_edn_arb.gen_normal_case.prio_mask_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_edn_arb.gen_normal_case.prio_mask_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_intr_esc0.intr_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_intr_esc0.intr_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_intr_esc1.intr_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_intr_esc1.intr_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.addr_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.addr_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.cnt_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.err_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.err_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.rdata_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.rdata_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.size_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.size_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_rdata_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_rdata_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_regfile_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_regfile_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_rvalid_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.tlul_rvalid_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.addr_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.addr_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rdata_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rdata_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.req_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.req_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rerror_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rerror_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rvalid_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rvalid_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rvalid_sram_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.rvalid_sram_q    &&
     //   top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.mem    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.mem &&
     //   top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.rdata_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.u_mem.gen_generic.u_impl_generic.rdata_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.wdata_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.wdata_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.wmask_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.wmask_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.write_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_prim_ram_1p_adv.write_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_state_regs.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_state_regs.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.intg_error_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.intg_error_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.valid_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.valid_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.wdata_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp.gen_generic.u_impl_generic.wdata_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_arb.gen_normal_case.prio_mask_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_arb.gen_normal_case.prio_mask_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_dai.base_sel_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_dai.base_sel_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_dai.cnt_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_dai.cnt_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_dai.data_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_dai.data_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_dai.error_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_dai.error_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_dai.u_state_regs.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_dai.u_state_regs.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.edn_req_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.edn_req_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.entropy_cnt_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.entropy_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.key_out_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.key_out_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.nonce_out_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.nonce_out_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.seed_cnt_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.seed_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.seed_valid_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.seed_valid_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.u_req_arb.gen_normal_case.prio_mask_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.u_req_arb.gen_normal_case.prio_mask_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_kdi.u_state_regs.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_kdi.u_state_regs.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lci.cnt_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lci.cnt_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lci.error_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lci.error_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lci.u_state_regs.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lci.u_state_regs.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.chk_timeout_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.chk_timeout_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.cnsty_chk_req_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.cnsty_chk_req_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.cnsty_chk_trig_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.cnsty_chk_trig_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[0].u_prim_flop_cnsty_cnt.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[0].u_prim_flop_cnsty_cnt.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[0].u_prim_flop_integ_cnt.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[0].u_prim_flop_integ_cnt.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[1].u_prim_flop_cnsty_cnt.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[1].u_prim_flop_cnsty_cnt.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[1].u_prim_flop_integ_cnt.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_cnt[1].u_prim_flop_integ_cnt.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.cnt_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.perturbed_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.gen_max_len_sva.perturbed_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.lfsr_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[0].u_prim_lfsr.lfsr_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.cnt_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.perturbed_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.gen_max_len_sva.perturbed_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.lfsr_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.gen_double_lfsr[1].u_prim_lfsr.lfsr_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.integ_chk_req_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.integ_chk_req_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.integ_chk_trig_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.integ_chk_trig_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.reseed_timer_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.reseed_timer_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_ctrl_lfsr_timer.u_state_regs.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_ctrl_lfsr_timer.u_state_regs.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_init_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_init_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_init_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_init_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_otp_rsp_fifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.fips_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.fips_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.clr_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.clr_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.data_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.data_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.depth_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_packer_fifo.depth_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_edn_req.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_check_byp_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_check_byp_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_check_byp_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_check_byp_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_creator_seed_sw_rw_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_creator_seed_sw_rw_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_creator_seed_sw_rw_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_creator_seed_sw_rw_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_dft_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_dft_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_dft_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_dft_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_escalate_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_seed_hw_rd_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_seed_hw_rd_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_prim_lc_sync_seed_hw_rd_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_prim_lc_sync_seed_hw_rd_en.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_regwen.q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_regwen.qe    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_timeout.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_timeout.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_timeout.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_timeout.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_trigger_regwen.q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_trigger_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_check_trigger_regwen.qe    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_check_trigger_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_consistency_check_period.q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_consistency_check_period.q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_consistency_check_period.qe    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_consistency_check_period.qe &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_creator_sw_cfg_read_lock.q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_creator_sw_cfg_read_lock.q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_creator_sw_cfg_read_lock.qe    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_creator_sw_cfg_read_lock.qe &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_address.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_address.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_address.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_address.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_wdata_0.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_wdata_0.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_wdata_0.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_wdata_0.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_wdata_1.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_wdata_1.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_direct_access_wdata_1.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_direct_access_wdata_1.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_integrity_check_period.q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_integrity_check_period.q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_integrity_check_period.qe  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_integrity_check_period.qe   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_enable_otp_error.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_enable_otp_error.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_enable_otp_error.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_enable_otp_error.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_enable_otp_operation_done.q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_enable_otp_operation_done.q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_enable_otp_operation_done.qe  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_enable_otp_operation_done.qe   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_state_otp_error.q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_state_otp_error.q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_state_otp_error.qe    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_state_otp_error.qe &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_state_otp_operation_done.q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_state_otp_operation_done.q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_intr_state_otp_operation_done.qe   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_intr_state_otp_operation_done.qe    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_owner_sw_cfg_read_lock.q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_owner_sw_cfg_read_lock.q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_owner_sw_cfg_read_lock.qe  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_owner_sw_cfg_read_lock.qe   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.dev_select_outstanding  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.dev_select_outstanding   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.err_resp.err_opcode == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.err_resp.err_opcode  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.err_resp.err_req_pending    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.err_resp.err_req_pending &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.err_resp.err_rsp_pending    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.err_resp.err_rsp_pending &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.err_resp.err_size   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.err_resp.err_size    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.err_resp.err_source == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.err_resp.err_source  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_reg.u_socket.num_req_outstanding == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_reg.u_socket.num_req_outstanding  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.cnt_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.cnt_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.data_shadow_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.data_shadow_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.data_state_q  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.data_state_q   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.digest_mode_q == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.digest_mode_q  &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.digest_state_q    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.digest_state_q &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.idx_state_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.idx_state_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.key_state_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.key_state_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.u_state_regs.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.u_state_regs.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl.valid_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl.valid_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_scrmbl_mtx.gen_normal_case.prio_mask_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_scrmbl_mtx.gen_normal_case.prio_mask_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.intg_error_q   == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.intg_error_q    &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_reqfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_rspfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_otp_ctrl.u_tlul_adapter_sram.u_sramreqfifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.alert_set_q == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.alert_set_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q    == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.ping_set_q  == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.ping_set_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.state_q == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.state_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q    == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q   == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o == top_level_upec.top_earlgrey_2.u_pattgen.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.bit_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.bit_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.clk_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.clk_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.complete_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.complete_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.complete_q2    == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.complete_q2 &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.data_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.data_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.len_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.len_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.pcl_int_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.pcl_int_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.polarity_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.polarity_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.prediv_q   == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.prediv_q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.rep_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.rep_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan0.reps_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan0.reps_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.bit_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.bit_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.clk_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.clk_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.complete_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.complete_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.complete_q2    == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.complete_q2 &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.data_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.data_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.len_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.len_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.pcl_int_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.pcl_int_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.polarity_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.polarity_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.prediv_q   == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.prediv_q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.rep_cnt_q  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.rep_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.chan1.reps_q == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.chan1.reps_q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.intr_hw_done_ch0.intr_o  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.intr_hw_done_ch0.intr_o   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_pattgen_core.intr_hw_done_ch1.intr_o  == top_level_upec.top_earlgrey_2.u_pattgen.u_pattgen_core.intr_hw_done_ch1.intr_o   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.intg_err_q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_enable_ch0.q   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_enable_ch0.q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_enable_ch0.qe  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_enable_ch0.qe   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_enable_ch1.q   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_enable_ch1.q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_enable_ch1.qe  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_enable_ch1.qe   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_polarity_ch0.q == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_polarity_ch0.q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_polarity_ch0.qe    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_polarity_ch0.qe &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_polarity_ch1.q == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_polarity_ch1.q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_ctrl_polarity_ch1.qe    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_ctrl_polarity_ch1.qe &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch0_0.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch0_0.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch0_0.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch0_0.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch0_1.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch0_1.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch0_1.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch0_1.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch1_0.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch1_0.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch1_0.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch1_0.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch1_1.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch1_1.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_data_ch1_1.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_data_ch1_1.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_enable_done_ch0.q  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_enable_done_ch0.q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_enable_done_ch0.qe == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_enable_done_ch0.qe  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_enable_done_ch1.q  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_enable_done_ch1.q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_enable_done_ch1.qe == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_enable_done_ch1.qe  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_state_done_ch0.q   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_state_done_ch0.q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_state_done_ch0.qe  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_state_done_ch0.qe   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_state_done_ch1.q   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_state_done_ch1.q    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_intr_state_done_ch1.qe  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_intr_state_done_ch1.qe   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_prediv_ch0.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_prediv_ch0.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_prediv_ch0.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_prediv_ch0.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_prediv_ch1.q    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_prediv_ch1.q &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_prediv_ch1.qe   == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_prediv_ch1.qe    &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_len_ch0.q  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_len_ch0.q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_len_ch0.qe == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_len_ch0.qe  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_len_ch1.q  == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_len_ch1.q   &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_len_ch1.qe == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_len_ch1.qe  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_reps_ch0.q == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_reps_ch0.q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_reps_ch0.qe    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_reps_ch0.qe &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_reps_ch1.q == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_reps_ch1.q  &&
        top_level_upec.top_earlgrey_1.u_pattgen.u_reg.u_size_reps_ch1.qe    == top_level_upec.top_earlgrey_2.u_pattgen.u_reg.u_size_reps_ch1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_oe_retreg_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_oe_retreg_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_out_retreg_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_out_retreg_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.dio_pad_attr_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.dio_pad_attr_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.alert_set_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.ping_set_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.state_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.state_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[0].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[1].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[2].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[3].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[4].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[5].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[6].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_cnt_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_filter_en_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_filter_en_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_filter_out_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_filter_out_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_cause_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_cause_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_cnt_th_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_cnt_th_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_mode_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.aon_wkup_mode_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_filter.stored_value_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_filter.stored_value_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_filter.stored_vector_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_filter.stored_vector_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_in.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_cause_out.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_flop_2sync_filter.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level   == top_level_upec.top_earlgrey_2.u_pinmux_aon.gen_wkup_detect[7].u_pinmux_wkup.i_prim_pulse_sync_cause.src_level    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_oe_retreg_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_oe_retreg_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_out_retreg_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_out_retreg_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.mio_pad_attr_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.mio_pad_attr_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.sleep_en_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.sleep_en_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.dft_strap_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.dft_strap_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.dft_strap_valid_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.dft_strap_valid_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.tap_strap_q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.tap_strap_q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_dft.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_dft.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_dft.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_dft.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_rv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_rv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_rv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_pinmux_strap_sampling.u_prim_lc_sync_rv.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_0.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_0.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_0.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_1.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_1.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_1.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_10.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_10.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_10.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_10.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_11.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_11.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_11.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_11.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_12.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_12.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_12.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_12.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_13.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_13.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_13.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_13.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_14.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_14.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_14.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_14.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_15.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_15.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_15.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_15.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_16.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_16.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_16.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_16.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_17.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_17.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_17.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_17.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_18.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_18.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_18.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_18.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_19.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_19.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_19.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_19.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_2.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_2.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_2.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_20.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_20.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_20.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_20.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_21.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_21.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_21.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_21.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_22.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_22.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_22.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_22.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_23.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_23.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_23.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_23.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_3.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_3.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_3.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_4.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_4.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_4.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_5.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_5.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_5.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_6.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_6.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_6.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_6.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_7.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_7.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_7.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_7.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_8.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_8.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_8.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_8.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_9.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_9.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_9.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_attr_regwen_9.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_10.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_10.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_10.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_10.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_11.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_11.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_11.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_11.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_12.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_12.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_12.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_12.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_13.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_13.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_13.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_13.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_14.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_14.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_14.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_14.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_15.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_15.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_15.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_15.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_16.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_16.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_16.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_16.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_17.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_17.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_17.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_17.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_18.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_18.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_18.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_18.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_19.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_19.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_19.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_19.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_20.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_20.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_20.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_20.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_21.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_21.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_21.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_21.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_22.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_22.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_22.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_22.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_23.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_23.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_23.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_23.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_8.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_8.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_8.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_8.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_9.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_9.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_9.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_en_9.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_0.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_0.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_0.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_1.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_1.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_1.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_10.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_10.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_10.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_10.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_11.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_11.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_11.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_11.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_12.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_12.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_12.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_12.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_13.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_13.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_13.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_13.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_14.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_14.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_14.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_14.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_15.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_15.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_15.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_15.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_16.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_16.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_16.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_16.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_17.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_17.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_17.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_17.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_18.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_18.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_18.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_18.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_19.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_19.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_19.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_19.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_2.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_2.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_2.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_20.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_20.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_20.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_20.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_21.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_21.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_21.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_21.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_22.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_22.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_22.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_22.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_23.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_23.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_23.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_23.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_3.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_3.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_3.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_4.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_4.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_4.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_5.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_5.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_5.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_6.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_6.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_6.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_6.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_7.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_7.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_7.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_7.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_8.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_8.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_8.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_8.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_9.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_9.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_9.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_mode_9.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_10.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_10.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_10.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_10.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_11.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_11.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_11.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_11.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_12.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_12.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_12.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_12.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_13.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_13.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_13.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_13.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_14.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_14.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_14.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_14.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_15.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_15.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_15.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_15.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_16.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_16.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_16.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_16.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_17.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_17.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_17.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_17.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_18.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_18.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_18.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_18.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_19.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_19.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_19.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_19.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_20.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_20.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_20.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_20.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_21.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_21.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_21.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_21.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_22.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_22.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_22.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_22.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_23.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_23.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_23.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_23.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_8.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_8.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_8.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_8.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_9.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_9.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_9.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_regwen_9.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_0.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_0.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_0.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_1.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_1.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_1.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_10.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_10.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_10.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_10.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_11.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_11.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_11.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_11.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_12.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_12.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_12.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_12.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_13.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_13.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_13.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_13.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_14.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_14.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_14.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_14.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_15.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_15.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_15.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_15.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_16.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_16.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_16.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_16.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_17.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_17.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_17.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_17.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_18.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_18.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_18.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_18.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_19.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_19.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_19.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_19.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_2.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_2.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_2.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_20.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_20.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_20.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_20.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_21.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_21.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_21.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_21.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_22.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_22.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_22.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_22.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_23.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_23.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_23.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_23.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_3.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_3.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_3.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_4.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_4.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_4.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_5.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_5.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_5.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_6.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_6.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_6.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_6.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_7.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_7.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_7.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_7.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_8.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_8.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_8.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_8.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_9.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_9.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_9.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_dio_pad_sleep_status_en_9.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_0.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_0.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_0.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_1.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_1.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_1.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_10.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_10.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_10.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_10.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_11.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_11.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_11.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_11.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_12.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_12.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_12.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_12.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_13.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_13.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_13.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_13.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_14.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_14.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_14.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_14.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_15.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_15.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_15.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_15.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_16.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_16.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_16.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_16.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_17.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_17.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_17.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_17.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_18.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_18.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_18.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_18.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_19.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_19.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_19.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_19.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_2.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_2.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_2.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_20.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_20.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_20.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_20.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_21.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_21.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_21.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_21.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_22.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_22.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_22.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_22.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_23.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_23.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_23.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_23.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_24.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_24.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_24.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_24.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_25.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_25.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_25.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_25.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_26.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_26.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_26.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_26.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_27.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_27.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_27.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_27.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_28.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_28.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_28.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_28.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_29.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_29.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_29.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_29.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_3.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_3.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_3.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_30.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_30.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_30.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_30.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_31.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_31.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_31.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_31.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_32.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_32.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_32.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_32.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_33.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_33.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_33.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_33.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_34.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_34.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_34.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_34.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_35.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_35.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_35.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_35.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_36.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_36.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_36.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_36.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_37.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_37.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_37.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_37.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_38.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_38.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_38.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_38.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_39.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_39.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_39.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_39.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_4.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_4.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_4.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_40.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_40.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_40.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_40.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_41.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_41.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_41.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_41.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_42.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_42.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_42.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_42.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_43.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_43.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_43.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_43.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_44.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_44.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_44.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_44.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_45.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_45.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_45.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_45.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_46.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_46.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_46.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_46.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_5.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_5.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_5.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_6.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_6.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_6.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_6.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_7.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_7.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_7.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_7.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_8.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_8.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_8.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_8.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_9.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_9.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_9.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_9.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_0.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_0.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_0.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_0.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_1.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_1.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_1.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_1.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_10.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_10.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_10.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_10.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_11.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_11.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_11.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_11.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_12.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_12.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_12.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_12.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_13.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_13.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_13.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_13.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_14.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_14.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_14.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_14.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_15.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_15.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_15.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_15.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_16.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_16.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_16.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_16.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_17.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_17.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_17.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_17.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_18.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_18.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_18.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_18.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_19.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_19.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_19.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_19.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_2.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_2.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_2.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_2.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_20.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_20.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_20.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_20.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_21.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_21.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_21.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_21.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_22.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_22.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_22.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_22.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_23.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_23.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_23.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_23.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_24.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_24.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_24.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_24.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_25.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_25.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_25.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_25.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_26.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_26.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_26.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_26.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_27.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_27.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_27.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_27.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_28.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_28.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_28.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_28.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_29.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_29.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_29.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_29.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_3.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_3.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_3.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_3.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_30.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_30.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_30.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_30.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_31.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_31.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_31.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_31.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_32.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_32.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_32.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_32.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_33.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_33.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_33.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_33.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_34.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_34.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_34.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_34.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_35.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_35.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_35.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_35.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_36.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_36.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_36.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_36.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_37.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_37.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_37.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_37.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_38.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_38.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_38.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_38.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_39.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_39.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_39.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_39.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_4.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_4.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_4.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_4.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_40.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_40.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_40.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_40.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_41.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_41.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_41.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_41.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_42.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_42.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_42.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_42.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_43.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_43.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_43.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_43.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_44.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_44.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_44.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_44.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_45.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_45.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_45.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_45.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_46.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_46.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_46.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_46.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_5.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_5.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_5.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_5.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_6.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_6.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_6.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_6.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_7.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_7.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_7.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_7.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_8.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_8.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_8.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_8.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_9.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_9.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_outsel_regwen_9.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_outsel_regwen_9.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_0.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_0.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_0.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_1.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_1.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_1.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_10.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_10.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_10.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_10.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_11.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_11.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_11.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_11.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_12.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_12.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_12.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_12.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_13.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_13.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_13.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_13.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_14.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_14.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_14.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_14.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_15.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_15.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_15.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_15.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_16.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_16.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_16.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_16.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_17.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_17.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_17.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_17.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_18.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_18.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_18.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_18.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_19.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_19.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_19.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_19.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_2.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_2.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_2.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_20.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_20.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_20.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_20.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_21.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_21.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_21.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_21.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_22.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_22.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_22.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_22.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_23.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_23.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_23.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_23.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_24.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_24.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_24.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_24.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_25.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_25.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_25.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_25.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_26.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_26.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_26.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_26.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_27.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_27.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_27.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_27.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_28.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_28.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_28.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_28.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_29.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_29.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_29.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_29.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_3.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_3.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_3.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_30.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_30.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_30.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_30.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_31.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_31.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_31.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_31.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_32.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_32.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_32.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_32.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_33.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_33.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_33.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_33.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_34.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_34.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_34.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_34.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_35.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_35.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_35.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_35.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_36.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_36.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_36.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_36.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_37.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_37.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_37.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_37.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_38.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_38.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_38.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_38.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_39.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_39.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_39.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_39.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_4.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_4.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_4.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_40.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_40.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_40.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_40.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_41.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_41.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_41.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_41.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_42.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_42.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_42.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_42.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_43.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_43.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_43.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_43.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_44.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_44.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_44.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_44.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_45.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_45.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_45.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_45.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_46.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_46.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_46.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_46.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_5.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_5.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_5.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_6.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_6.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_6.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_6.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_7.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_7.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_7.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_7.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_8.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_8.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_8.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_8.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_9.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_9.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_9.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_attr_regwen_9.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_10.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_10.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_10.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_10.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_11.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_11.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_11.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_11.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_12.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_12.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_12.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_12.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_13.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_13.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_13.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_13.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_14.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_14.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_14.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_14.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_15.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_15.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_15.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_15.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_16.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_16.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_16.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_16.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_17.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_17.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_17.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_17.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_18.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_18.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_18.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_18.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_19.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_19.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_19.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_19.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_20.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_20.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_20.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_20.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_21.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_21.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_21.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_21.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_22.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_22.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_22.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_22.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_23.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_23.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_23.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_23.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_24.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_24.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_24.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_24.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_25.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_25.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_25.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_25.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_26.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_26.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_26.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_26.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_27.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_27.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_27.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_27.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_28.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_28.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_28.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_28.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_29.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_29.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_29.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_29.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_30.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_30.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_30.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_30.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_31.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_31.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_31.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_31.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_32.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_32.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_32.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_32.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_33.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_33.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_33.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_33.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_34.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_34.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_34.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_34.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_35.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_35.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_35.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_35.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_36.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_36.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_36.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_36.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_37.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_37.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_37.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_37.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_38.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_38.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_38.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_38.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_39.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_39.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_39.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_39.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_40.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_40.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_40.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_40.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_41.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_41.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_41.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_41.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_42.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_42.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_42.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_42.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_43.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_43.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_43.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_43.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_44.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_44.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_44.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_44.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_45.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_45.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_45.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_45.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_46.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_46.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_46.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_46.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_8.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_8.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_8.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_8.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_9.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_9.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_9.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_en_9.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_0.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_0.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_0.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_1.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_1.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_1.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_10.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_10.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_10.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_10.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_11.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_11.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_11.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_11.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_12.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_12.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_12.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_12.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_13.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_13.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_13.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_13.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_14.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_14.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_14.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_14.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_15.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_15.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_15.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_15.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_16.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_16.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_16.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_16.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_17.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_17.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_17.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_17.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_18.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_18.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_18.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_18.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_19.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_19.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_19.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_19.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_2.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_2.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_2.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_20.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_20.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_20.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_20.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_21.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_21.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_21.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_21.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_22.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_22.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_22.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_22.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_23.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_23.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_23.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_23.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_24.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_24.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_24.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_24.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_25.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_25.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_25.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_25.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_26.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_26.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_26.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_26.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_27.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_27.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_27.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_27.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_28.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_28.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_28.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_28.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_29.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_29.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_29.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_29.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_3.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_3.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_3.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_30.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_30.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_30.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_30.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_31.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_31.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_31.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_31.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_32.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_32.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_32.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_32.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_33.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_33.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_33.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_33.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_34.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_34.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_34.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_34.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_35.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_35.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_35.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_35.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_36.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_36.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_36.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_36.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_37.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_37.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_37.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_37.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_38.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_38.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_38.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_38.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_39.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_39.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_39.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_39.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_4.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_4.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_4.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_40.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_40.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_40.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_40.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_41.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_41.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_41.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_41.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_42.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_42.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_42.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_42.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_43.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_43.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_43.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_43.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_44.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_44.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_44.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_44.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_45.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_45.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_45.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_45.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_46.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_46.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_46.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_46.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_5.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_5.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_5.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_6.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_6.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_6.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_6.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_7.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_7.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_7.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_7.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_8.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_8.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_8.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_8.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_9.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_9.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_9.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_mode_9.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_10.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_10.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_10.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_10.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_11.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_11.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_11.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_11.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_12.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_12.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_12.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_12.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_13.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_13.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_13.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_13.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_14.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_14.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_14.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_14.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_15.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_15.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_15.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_15.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_16.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_16.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_16.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_16.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_17.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_17.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_17.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_17.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_18.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_18.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_18.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_18.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_19.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_19.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_19.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_19.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_20.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_20.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_20.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_20.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_21.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_21.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_21.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_21.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_22.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_22.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_22.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_22.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_23.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_23.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_23.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_23.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_24.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_24.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_24.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_24.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_25.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_25.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_25.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_25.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_26.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_26.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_26.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_26.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_27.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_27.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_27.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_27.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_28.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_28.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_28.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_28.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_29.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_29.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_29.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_29.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_30.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_30.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_30.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_30.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_31.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_31.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_31.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_31.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_32.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_32.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_32.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_32.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_33.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_33.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_33.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_33.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_34.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_34.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_34.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_34.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_35.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_35.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_35.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_35.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_36.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_36.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_36.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_36.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_37.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_37.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_37.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_37.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_38.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_38.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_38.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_38.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_39.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_39.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_39.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_39.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_40.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_40.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_40.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_40.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_41.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_41.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_41.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_41.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_42.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_42.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_42.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_42.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_43.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_43.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_43.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_43.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_44.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_44.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_44.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_44.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_45.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_45.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_45.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_45.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_46.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_46.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_46.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_46.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_8.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_8.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_8.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_8.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_9.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_9.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_9.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_regwen_9.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_0.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_0.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_0.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_0.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_1.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_1.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_1.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_1.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_10.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_10.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_10.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_10.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_11.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_11.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_11.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_11.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_12.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_12.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_12.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_12.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_13.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_13.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_13.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_13.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_14.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_14.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_14.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_14.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_15.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_15.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_15.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_15.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_16.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_16.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_16.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_16.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_17.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_17.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_17.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_17.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_18.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_18.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_18.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_18.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_19.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_19.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_19.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_19.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_2.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_2.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_2.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_2.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_20.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_20.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_20.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_20.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_21.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_21.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_21.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_21.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_22.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_22.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_22.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_22.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_23.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_23.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_23.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_23.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_24.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_24.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_24.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_24.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_25.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_25.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_25.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_25.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_26.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_26.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_26.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_26.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_27.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_27.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_27.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_27.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_28.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_28.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_28.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_28.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_29.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_29.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_29.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_29.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_3.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_3.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_3.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_3.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_30.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_30.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_30.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_30.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_31.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_31.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_31.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_31.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_4.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_4.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_4.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_4.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_5.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_5.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_5.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_5.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_6.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_6.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_6.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_6.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_7.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_7.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_7.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_7.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_8.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_8.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_8.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_8.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_9.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_9.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_9.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_0_en_9.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_32.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_32.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_32.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_32.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_33.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_33.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_33.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_33.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_34.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_34.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_34.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_34.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_35.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_35.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_35.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_35.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_36.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_36.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_36.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_36.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_37.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_37.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_37.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_37.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_38.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_38.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_38.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_38.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_39.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_39.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_39.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_39.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_40.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_40.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_40.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_40.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_41.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_41.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_41.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_41.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_42.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_42.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_42.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_42.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_43.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_43.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_43.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_43.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_44.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_44.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_44.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_44.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_45.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_45.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_45.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_45.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_46.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_46.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_46.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_pad_sleep_status_1_en_46.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_10.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_10.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_10.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_10.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_11.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_11.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_11.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_11.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_12.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_12.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_12.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_12.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_13.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_13.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_13.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_13.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_14.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_14.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_14.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_14.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_15.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_15.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_15.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_15.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_16.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_16.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_16.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_16.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_17.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_17.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_17.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_17.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_18.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_18.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_18.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_18.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_19.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_19.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_19.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_19.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_20.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_20.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_20.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_20.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_21.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_21.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_21.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_21.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_22.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_22.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_22.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_22.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_23.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_23.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_23.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_23.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_24.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_24.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_24.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_24.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_25.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_25.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_25.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_25.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_26.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_26.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_26.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_26.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_27.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_27.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_27.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_27.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_28.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_28.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_28.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_28.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_29.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_29.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_29.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_29.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_30.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_30.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_30.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_30.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_31.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_31.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_31.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_31.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_32.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_32.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_32.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_32.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_33.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_33.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_33.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_33.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_34.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_34.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_34.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_34.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_35.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_35.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_35.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_35.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_36.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_36.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_36.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_36.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_37.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_37.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_37.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_37.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_38.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_38.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_38.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_38.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_39.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_39.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_39.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_39.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_40.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_40.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_40.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_40.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_41.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_41.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_41.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_41.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_42.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_42.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_42.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_42.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_43.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_43.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_43.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_43.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_44.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_44.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_44.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_44.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_45.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_45.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_45.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_45.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_46.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_46.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_46.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_46.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_47.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_47.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_47.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_47.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_48.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_48.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_48.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_48.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_49.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_49.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_49.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_49.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_50.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_50.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_50.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_50.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_51.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_51.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_51.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_51.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_52.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_52.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_52.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_52.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_53.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_53.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_53.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_53.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_54.q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_54.q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_54.qe   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_54.qe    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_8.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_8.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_8.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_8.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_9.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_9.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_9.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_9.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_0.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_0.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_0.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_1.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_1.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_1.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_10.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_10.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_10.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_10.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_11.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_11.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_11.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_11.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_12.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_12.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_12.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_12.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_13.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_13.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_13.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_13.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_14.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_14.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_14.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_14.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_15.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_15.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_15.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_15.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_16.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_16.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_16.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_16.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_17.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_17.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_17.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_17.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_18.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_18.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_18.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_18.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_19.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_19.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_19.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_19.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_2.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_2.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_2.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_20.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_20.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_20.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_20.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_21.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_21.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_21.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_21.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_22.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_22.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_22.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_22.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_23.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_23.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_23.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_23.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_24.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_24.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_24.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_24.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_25.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_25.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_25.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_25.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_26.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_26.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_26.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_26.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_27.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_27.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_27.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_27.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_28.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_28.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_28.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_28.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_29.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_29.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_29.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_29.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_3.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_3.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_3.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_30.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_30.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_30.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_30.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_31.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_31.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_31.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_31.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_32.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_32.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_32.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_32.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_33.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_33.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_33.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_33.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_34.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_34.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_34.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_34.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_35.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_35.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_35.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_35.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_36.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_36.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_36.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_36.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_37.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_37.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_37.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_37.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_38.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_38.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_38.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_38.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_39.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_39.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_39.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_39.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_4.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_4.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_4.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_40.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_40.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_40.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_40.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_41.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_41.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_41.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_41.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_42.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_42.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_42.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_42.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_43.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_43.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_43.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_43.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_44.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_44.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_44.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_44.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_45.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_45.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_45.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_45.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_46.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_46.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_46.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_46.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_47.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_47.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_47.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_47.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_48.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_48.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_48.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_48.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_49.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_49.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_49.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_49.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_5.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_5.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_5.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_50.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_50.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_50.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_50.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_51.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_51.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_51.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_51.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_52.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_52.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_52.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_52.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_53.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_53.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_53.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_53.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_54.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_54.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_54.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_54.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_6.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_6.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_6.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_6.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_7.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_7.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_7.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_7.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_8.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_8.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_8.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_8.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_9.q  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_9.q   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_9.qe == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_mio_periph_insel_regwen_9.qe  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_filter_0.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_filter_0.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_filter_0.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_filter_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_miodio_0.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_miodio_0.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_miodio_0.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_miodio_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_mode_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_mode_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_0_mode_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_0_mode_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_filter_1.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_filter_1.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_filter_1.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_filter_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_miodio_1.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_miodio_1.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_miodio_1.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_miodio_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_mode_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_mode_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_1_mode_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_1_mode_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_filter_2.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_filter_2.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_filter_2.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_filter_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_miodio_2.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_miodio_2.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_miodio_2.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_miodio_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_mode_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_mode_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_2_mode_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_2_mode_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_filter_3.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_filter_3.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_filter_3.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_filter_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_miodio_3.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_miodio_3.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_miodio_3.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_miodio_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_mode_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_mode_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_3_mode_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_3_mode_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_filter_4.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_filter_4.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_filter_4.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_filter_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_miodio_4.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_miodio_4.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_miodio_4.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_miodio_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_mode_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_mode_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_4_mode_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_4_mode_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_filter_5.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_filter_5.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_filter_5.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_filter_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_miodio_5.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_miodio_5.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_miodio_5.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_miodio_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_mode_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_mode_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_5_mode_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_5_mode_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_filter_6.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_filter_6.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_filter_6.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_filter_6.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_miodio_6.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_miodio_6.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_miodio_6.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_miodio_6.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_mode_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_mode_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_6_mode_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_6_mode_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_filter_7.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_filter_7.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_filter_7.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_filter_7.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_miodio_7.q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_miodio_7.q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_miodio_7.qe  == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_miodio_7.qe   &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_mode_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_mode_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_7_mode_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_7_mode_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_cnt_th_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_en_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_en_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_padsel_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_padsel_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_0.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_0.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_0.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_0.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_1.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_1.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_1.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_1.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_2.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_2.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_2.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_2.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_3.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_3.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_3.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_3.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_4.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_4.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_4.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_4.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_5.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_5.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_5.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_5.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_6.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_6.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_6.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_6.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_7.q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_7.q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_reg.u_wkup_detector_regwen_7.qe    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_reg.u_wkup_detector_regwen_7.qe &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.astate_q   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.astate_q    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.filter_activity.stored_value_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.filter_activity.stored_value_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.filter_activity.stored_vector_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.filter_activity.stored_vector_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[0].u_filter.stored_value_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[0].u_filter.stored_value_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[0].u_filter.stored_vector_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[0].u_filter.stored_vector_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[1].u_filter.stored_value_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[1].u_filter.stored_value_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[1].u_filter.stored_vector_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[1].u_filter.stored_vector_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[2].u_filter.stored_value_q == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[2].u_filter.stored_value_q  &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[2].u_filter.stored_vector_q    == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.gen_filters[2].u_filter.stored_vector_q &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.u_cdc_suspend_req.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.u_cdc_suspend_req.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pinmux_aon.u_usbdev_aon_wake.u_cdc_suspend_req.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pinmux_aon.u_usbdev_aon_wake.u_cdc_suspend_req.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.beat_ctr_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.beat_ctr_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[0].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[1].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[2].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[3].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[4].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.blink_ctr_q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.blink_ctr_q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.dc_htbt_q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.dc_htbt_q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.htbt_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.htbt_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.htbt_direction  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.gen_chan_insts[5].u_chan.htbt_direction   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.phase_ctr_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.phase_ctr_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.common_sync_q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.common_sync_q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[0].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[1].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[2].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[3].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[4].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].chan_sync_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].chan_sync_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].u_common_sync2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.gen_chan_cdc[5].u_common_sync2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.u_common_sync1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.u_common_sync1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_pwm_core.u_pwm_cdc.u_common_sync1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_pwm_core.u_pwm_cdc.u_common_sync1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.intg_err_q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_0_x_0.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_0_x_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_0_x_0.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_0_x_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_0_y_0.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_0_y_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_0_y_0.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_0_y_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_1_x_1.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_1_x_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_1_x_1.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_1_x_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_1_y_1.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_1_y_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_1_y_1.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_1_y_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_2_x_2.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_2_x_2.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_2_x_2.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_2_x_2.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_2_y_2.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_2_y_2.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_2_y_2.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_2_y_2.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_3_x_3.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_3_x_3.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_3_x_3.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_3_x_3.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_3_y_3.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_3_y_3.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_3_y_3.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_3_y_3.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_4_x_4.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_4_x_4.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_4_x_4.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_4_x_4.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_4_y_4.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_4_y_4.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_4_y_4.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_4_y_4.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_5_x_5.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_5_x_5.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_5_x_5.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_5_x_5.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_5_y_5.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_5_y_5.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_blink_param_5_y_5.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_blink_param_5_y_5.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_clk_div.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_clk_div.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_clk_div.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_clk_div.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_cntr_en.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_cntr_en.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_cntr_en.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_cntr_en.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_dc_resn.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_dc_resn.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_cfg_dc_resn.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_cfg_dc_resn.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_0_a_0.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_0_a_0.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_0_a_0.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_0_a_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_0_b_0.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_0_b_0.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_0_b_0.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_0_b_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_1_a_1.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_1_a_1.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_1_a_1.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_1_a_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_1_b_1.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_1_b_1.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_1_b_1.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_1_b_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_2_a_2.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_2_a_2.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_2_a_2.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_2_a_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_2_b_2.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_2_b_2.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_2_b_2.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_2_b_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_3_a_3.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_3_a_3.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_3_a_3.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_3_a_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_3_b_3.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_3_b_3.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_3_b_3.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_3_b_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_4_a_4.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_4_a_4.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_4_a_4.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_4_a_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_4_b_4.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_4_b_4.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_4_b_4.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_4_b_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_5_a_5.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_5_a_5.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_5_a_5.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_5_a_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_5_b_5.q  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_5_b_5.q   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_duty_cycle_5_b_5.qe == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_duty_cycle_5_b_5.qe  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_0.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_0.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_0.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_1.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_1.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_1.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_2.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_2.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_2.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_3.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_3.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_3.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_4.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_4.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_4.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_5.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_5.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_invert_invert_5.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_invert_invert_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_0.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_0.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_0.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_0.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_1.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_1.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_1.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_1.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_2.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_2.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_2.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_2.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_3.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_3.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_3.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_3.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_4.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_4.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_4.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_4.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_5.q   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_5.q    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_en_en_5.qe  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_en_en_5.qe   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_blink_en_0.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_blink_en_0.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_blink_en_0.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_blink_en_0.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_htbt_en_0.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_htbt_en_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_htbt_en_0.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_htbt_en_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_phase_delay_0.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_phase_delay_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_0_phase_delay_0.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_0_phase_delay_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_blink_en_1.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_blink_en_1.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_blink_en_1.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_blink_en_1.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_htbt_en_1.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_htbt_en_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_htbt_en_1.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_htbt_en_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_phase_delay_1.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_phase_delay_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_1_phase_delay_1.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_1_phase_delay_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_blink_en_2.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_blink_en_2.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_blink_en_2.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_blink_en_2.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_htbt_en_2.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_htbt_en_2.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_htbt_en_2.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_htbt_en_2.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_phase_delay_2.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_phase_delay_2.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_2_phase_delay_2.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_2_phase_delay_2.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_blink_en_3.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_blink_en_3.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_blink_en_3.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_blink_en_3.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_htbt_en_3.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_htbt_en_3.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_htbt_en_3.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_htbt_en_3.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_phase_delay_3.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_phase_delay_3.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_3_phase_delay_3.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_3_phase_delay_3.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_blink_en_4.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_blink_en_4.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_blink_en_4.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_blink_en_4.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_htbt_en_4.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_htbt_en_4.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_htbt_en_4.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_htbt_en_4.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_phase_delay_4.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_phase_delay_4.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_4_phase_delay_4.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_4_phase_delay_4.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_blink_en_5.q    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_blink_en_5.q &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_blink_en_5.qe   == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_blink_en_5.qe    &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_htbt_en_5.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_htbt_en_5.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_htbt_en_5.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_htbt_en_5.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_phase_delay_5.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_phase_delay_5.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_pwm_param_5_phase_delay_5.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_pwm_param_5_phase_delay_5.qe &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_regen.q == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_regen.q  &&
        top_level_upec.top_earlgrey_1.u_pwm_aon.u_reg.u_regen.qe    == top_level_upec.top_earlgrey_2.u_pwm_aon.u_reg.u_regen.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ack_pwrdn_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ack_pwrdn_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ack_pwrdn_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ack_pwrdn_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ack_pwrup_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ack_pwrup_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ack_pwrup_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ack_pwrup_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ast_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ast_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ast_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ast_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ext_req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ext_req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_ext_req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_ext_req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_pwrup_chg_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_pwrup_chg_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_pwrup_chg_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_pwrup_chg_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_req_pwrdn_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_req_pwrdn_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_req_pwrdn_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_req_pwrdn_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_req_pwrup_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_req_pwrup_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_req_pwrup_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_req_pwrup_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_scdc_sync.dst_level_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_scdc_sync.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_scdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_scdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_scdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_scdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_scdc_sync.src_level  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_scdc_sync.src_level   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.dst_level_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.src_level  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_cdc_sync.src_level   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_ext_req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_ext_req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.i_slow_ext_req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.i_slow_ext_req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.pwrup_cause_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.pwrup_cause_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.pwrup_cause_toggle_q2  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.pwrup_cause_toggle_q2   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_ast_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_ast_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_ast_q2    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_ast_q2 &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_core_clk_en_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_core_clk_en_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_io_clk_en_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_io_clk_en_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_main_pd_no    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_main_pd_no &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_reset_en_o    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_reset_en_o &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_usb_clk_en_active_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_usb_clk_en_active_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_usb_clk_en_lp_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_usb_clk_en_lp_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.slow_wakeup_en_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.slow_wakeup_en_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_flash_idle.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_flash_idle.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_flash_idle.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_flash_idle.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_otp.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_otp.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_otp.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_otp.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_rom_ctrl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_rom_ctrl.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_cdc.u_sync_rom_ctrl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_cdc.u_sync_rom_ctrl.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.ack_pwrup_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.ack_pwrup_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.ip_clk_en_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.ip_clk_en_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.low_power_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.low_power_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.req_pwrdn_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.req_pwrdn_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.reset_cause_q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.reset_cause_q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.reset_ongoing_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.reset_ongoing_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.rst_lc_req_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.rst_lc_req_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.rst_sys_req_q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.rst_sys_req_q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.state_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.state_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.strap_sampled  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.strap_sampled   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_fetch_en.u_prim_flop.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_fetch_en.u_prim_flop.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_reg_lc_init.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_reg_lc_init.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_reg_otp_init.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_reg_otp_init.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_slow_sync_lc_done.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_slow_sync_lc_done.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_slow_sync_lc_done.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_slow_sync_lc_done.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_sync_lc_done.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_sync_lc_done.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_fsm.u_sync_lc_done.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_fsm.u_sync_lc_done.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.ack_pwrdn_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.ack_pwrdn_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.cause_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.cause_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.cause_toggle_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.cause_toggle_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.core_clk_en_q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.core_clk_en_q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.io_clk_en_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.io_clk_en_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.pd_nq == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.pd_nq  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.pwr_clamp_env_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.pwr_clamp_env_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.pwr_clamp_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.pwr_clamp_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.req_pwrup_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.req_pwrup_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.state_q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.state_q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_slow_fsm.usb_clk_en_q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_slow_fsm.usb_clk_en_q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_wake_info.info == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_wake_info.info  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_wake_info.record_en    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_wake_info.record_en &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.i_wake_info.start_capture_q1 == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.i_wake_info.start_capture_q1  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.intr_wakeup.intr_o   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.intr_wakeup.intr_o    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.lowpwr_cfg_wen   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.lowpwr_cfg_wen    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_esc_rx.state_q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_esc_rx.state_q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_esc_rx.u_decode_esc.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_esc_rx.u_decode_esc.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_esc_rx.u_decode_esc.level_q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_esc_rx.u_decode_esc.level_q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_esc_rx.u_prim_generic_flop.q_o == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_esc_rx.u_prim_generic_flop.q_o  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_cfg_cdc_sync.q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_cfg_cdc_sync.q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_cfg_cdc_sync.qe  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_cfg_cdc_sync.qe   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_core_clk_en.q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_core_clk_en.q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_core_clk_en.qe   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_core_clk_en.qe    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_io_clk_en.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_io_clk_en.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_io_clk_en.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_io_clk_en.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_low_power_hint.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_low_power_hint.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_low_power_hint.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_low_power_hint.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_main_pd_n.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_main_pd_n.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_main_pd_n.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_main_pd_n.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_active.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_active.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_active.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_active.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_lp.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_lp.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_lp.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_control_usb_clk_en_lp.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_escalate_reset_status.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_escalate_reset_status.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_escalate_reset_status.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_escalate_reset_status.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_intr_enable.q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_intr_enable.q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_intr_enable.qe   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_intr_enable.qe    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_intr_state.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_intr_state.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_intr_state.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_intr_state.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_en_0.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_en_0.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_en_0.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_en_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_en_1.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_en_1.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_en_1.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_en_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_regwen.q    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_regwen.q &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_en_regwen.qe   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_en_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_status_val_0.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_status_val_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_status_val_0.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_status_val_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_status_val_1.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_status_val_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_reset_status_val_1.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_reset_status_val_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_info_capture_dis.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_info_capture_dis.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_info_capture_dis.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_info_capture_dis.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_0.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_0.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_0.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_0.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_1.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_1.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_1.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_1.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_2.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_2.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_2.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_2.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_3.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_3.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_3.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_3.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_4.q  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_4.q   &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wake_status_val_4.qe == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wake_status_val_4.qe  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_0.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_0.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_0.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_0.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_1.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_1.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_1.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_1.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_2.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_2.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_2.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_2.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_3.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_3.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_3.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_3.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_4.q == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_4.q  &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_en_4.qe    == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_en_4.qe &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_regwen.q   == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_regwen.q    &&
        top_level_upec.top_earlgrey_1.u_pwrmgr_aon.u_reg.u_wakeup_en_regwen.qe  == top_level_upec.top_earlgrey_2.u_pwrmgr_aon.u_reg.u_wakeup_en_regwen.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.first_reset  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.first_reset   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.cnt  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.cnt   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_filter_n == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_filter_n  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.rst_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.u_rst_flop.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_rst_por_aon[0].gen_rst_por_aon_normal.u_rst_por_aon.u_rst_flop.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[0].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[0].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[0].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[0].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[1].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[1].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[1].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[1].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[2].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[2].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[2].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[2].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[3].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[3].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[3].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[3].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[4].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[4].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[4].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[4].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[5].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[5].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[5].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[5].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[6].u_rst_sw_ctrl_reg.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[6].u_rst_sw_ctrl_reg.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.gen_sw_rst_ext_regs[6].u_rst_sw_ctrl_reg.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.gen_sw_rst_ext_regs[6].u_rst_sw_ctrl_reg.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_i2c2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_i2c2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_lc_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_lc_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_lc_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_lc_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_device.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_device.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_device.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_device.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_host0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_host0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_host0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_host0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_host1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_host1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_spi_host1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_spi_host1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys_aon.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys_aon.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys_aon.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys_aon.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_sys_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_sys_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_0_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_0_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_alert_info.slots_q == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_alert_info.slots_q  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io_div2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io_div2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io_div2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io_div2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_por_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_por_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_sys_aon.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_sys_aon.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_sys_aon.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_sys_aon.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_sys_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_sys_io_div4.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_aon_sys_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_aon_sys_io_div4.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_cpu_info.slots_q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_cpu_info.slots_q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_cpu_reset_synced.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_cpu_reset_synced.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_cpu_reset_synced.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_cpu_reset_synced.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_lc_src.gen_rst_pd_n[0].u_pd_rst.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_lc_src.gen_rst_pd_n[0].u_pd_rst.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_lc_src.u_aon_rst.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_lc_src.u_aon_rst.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_lc_src.u_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_lc_src.u_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_lc_src.u_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_lc_src.u_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_info_ctrl_en.q == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_info_ctrl_en.q  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_info_ctrl_en.qe    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_info_ctrl_en.qe &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_info_ctrl_index.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_info_ctrl_index.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_info_ctrl_index.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_info_ctrl_index.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_regwen.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_regwen.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_alert_regwen.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_alert_regwen.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_en.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_en.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_en.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_en.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_index.q    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_index.q &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_index.qe   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_info_ctrl_index.qe    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_regwen.q == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_cpu_regwen.qe    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_cpu_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_hw_req.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_hw_req.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_hw_req.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_hw_req.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_low_power_exit.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_low_power_exit.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_low_power_exit.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_low_power_exit.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_ndm_reset.q   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_ndm_reset.q    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_ndm_reset.qe  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_ndm_reset.qe   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_por.q == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_por.q  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_reset_info_por.qe    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_reset_info_por.qe &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_0.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_0.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_0.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_0.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_1.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_1.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_1.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_1.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_2.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_2.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_2.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_2.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_3.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_3.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_3.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_3.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_4.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_4.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_4.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_4.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_5.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_5.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_5.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_5.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_6.q  == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_6.q   &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_6.qe == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_reg.u_sw_rst_regen_en_6.qe  &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sys_src.gen_rst_pd_n[0].u_pd_rst.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sys_src.gen_rst_pd_n[0].u_pd_rst.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sys_src.u_aon_rst.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sys_src.u_aon_rst.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sys_src.u_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sys_src.u_lc.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rstmgr_aon.u_sys_src.u_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_rstmgr_aon.u_sys_src.u_lc.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_rv_timer.gen_harts[0].u_core.tick_count == top_level_upec.top_earlgrey_2.u_rv_timer.gen_harts[0].u_core.tick_count  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.gen_harts[0].u_intr_hw.intr_o  == top_level_upec.top_earlgrey_2.u_rv_timer.gen_harts[0].u_intr_hw.intr_o   &&
        top_level_upec.top_earlgrey_1.u_rv_timer.gen_harts[1].u_core.tick_count == top_level_upec.top_earlgrey_2.u_rv_timer.gen_harts[1].u_core.tick_count  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.gen_harts[1].u_intr_hw.intr_o  == top_level_upec.top_earlgrey_2.u_rv_timer.gen_harts[1].u_intr_hw.intr_o   &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.intg_err_q   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.intg_err_q    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_cfg0_prescale.q    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_cfg0_prescale.q &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_cfg0_prescale.qe   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_cfg0_prescale.qe    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_cfg0_step.q    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_cfg0_step.q &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_cfg0_step.qe   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_cfg0_step.qe    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_compare_lower0_0.q == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_compare_lower0_0.q  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_compare_lower0_0.qe    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_compare_lower0_0.qe &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_compare_upper0_0.q == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_compare_upper0_0.q  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_compare_upper0_0.qe    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_compare_upper0_0.qe &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_ctrl.q == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_ctrl.q  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_ctrl.qe    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_ctrl.qe &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_intr_enable0.q == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_intr_enable0.q  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_intr_enable0.qe    == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_intr_enable0.qe &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_intr_state0.q  == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_intr_state0.q   &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_intr_state0.qe == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_intr_state0.qe  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.error   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.error    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.outstanding == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.outstanding  &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.rdata   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.rdata    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.reqid   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.reqid    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.reqsz   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.reqsz    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_reg_if.rspop   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_reg_if.rspop    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_timer_v_lower0.q   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_timer_v_lower0.q    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_timer_v_lower0.qe  == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_timer_v_lower0.qe   &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_timer_v_upper0.q   == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_timer_v_upper0.q    &&
        top_level_upec.top_earlgrey_1.u_rv_timer.u_reg.u_timer_v_upper0.qe  == top_level_upec.top_earlgrey_2.u_rv_timer.u_reg.u_timer_v_upper0.qe   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[0].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[10].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[1].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[2].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[3].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[4].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[5].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[6].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[7].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[8].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.alert_set_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.alert_set_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.alert_test_set_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.alert_test_set_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.ping_set_q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.ping_set_q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.state_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.state_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ack.level_q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ack.level_q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ping.level_q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_decode_ping.level_q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_prim_generic_flop.q_o    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.gen_alert_senders[9].u_prim_alert_sender.u_prim_generic_flop.q_o &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.intg_err_q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_0.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_0.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_0.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_1.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_1.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_1.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_10.q   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_10.q    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_10.qe  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_10.qe   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_2.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_2.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_2.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_2.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_3.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_3.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_3.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_3.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_4.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_4.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_4.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_4.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_5.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_5.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_5.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_5.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_6.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_6.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_6.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_6.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_7.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_7.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_7.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_7.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_8.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_8.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_8.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_8.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_9.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_9.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_9.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_ack_mode_val_9.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_0.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_0.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_0.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_0.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_1.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_1.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_1.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_1.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_10.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_10.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_10.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_10.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_2.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_2.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_2.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_2.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_3.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_3.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_3.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_3.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_4.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_4.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_4.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_4.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_5.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_5.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_5.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_5.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_6.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_6.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_6.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_6.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_7.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_7.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_7.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_7.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_8.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_8.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_8.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_8.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_9.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_9.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_state_val_9.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_state_val_9.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_0.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_0.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_0.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_0.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_1.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_1.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_1.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_1.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_10.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_10.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_10.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_10.qe &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_2.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_2.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_2.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_2.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_3.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_3.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_3.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_3.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_4.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_4.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_4.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_4.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_5.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_5.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_5.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_5.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_6.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_6.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_6.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_6.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_7.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_7.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_7.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_7.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_8.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_8.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_8.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_8.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_9.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_9.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_9.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_alert_trig_val_9.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_cfg_regwen.q    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_cfg_regwen.q &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_cfg_regwen.qe   == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_cfg_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_status_ast_init_done.q  == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_status_ast_init_done.q   &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_status_ast_init_done.qe == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_status_ast_init_done.qe  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_status_io_pok.q == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_status_io_pok.q  &&
        top_level_upec.top_earlgrey_1.u_sensor_ctrl_aon.u_reg.u_status_io_pok.qe    == top_level_upec.top_earlgrey_2.u_sensor_ctrl_aon.u_reg.u_status_io_pok.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.cmd_dp_sel_outclk    == top_level_upec.top_earlgrey_2.u_spi_device.cmd_dp_sel_outclk &&
        top_level_upec.top_earlgrey_1.u_spi_device.fwm_rxerr_q  == top_level_upec.top_earlgrey_2.u_spi_device.fwm_rxerr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.alert_set_q  == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.ping_set_q   == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.state_q  == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.state_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q    == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q &&
        top_level_upec.top_earlgrey_1.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.io_mode_outclk   == top_level_upec.top_earlgrey_2.u_spi_device.io_mode_outclk    &&
        top_level_upec.top_earlgrey_1.u_spi_device.rxf_full_q   == top_level_upec.top_earlgrey_2.u_spi_device.rxf_full_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.rxlvl    == top_level_upec.top_earlgrey_2.u_spi_device.rxlvl &&
        top_level_upec.top_earlgrey_1.u_spi_device.sram_rxf_full_q  == top_level_upec.top_earlgrey_2.u_spi_device.sram_rxf_full_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.txf_empty_q  == top_level_upec.top_earlgrey_2.u_spi_device.txf_empty_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.txlvl    == top_level_upec.top_earlgrey_2.u_spi_device.txlvl &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_cmdparse.opcode_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_cmdparse.opcode_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_cmdparse.st    == top_level_upec.top_earlgrey_2.u_spi_device.u_cmdparse.st &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_fwmode_arb.gen_arb_ppc.u_reqarb.gen_normal_case.mask  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_fwmode_arb.gen_arb_ppc.u_reqarb.gen_normal_case.mask   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_fwmode_arb.u_req_fifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_gray_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_sync_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.fifo_rptr_sync_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.fifo_wptr_gray_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.fifo_wptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.fifo_wptr_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.fifo_wptr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.storage   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.byte_enable  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.byte_enable   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.cur_timer    == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.cur_timer &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.pos  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.pos   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.sram_req == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.sram_req  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.sram_wdata   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.sram_wdata    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.sram_write   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.sram_write    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.st   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.st    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_rxf_ctrl.wptr == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_rxf_ctrl.wptr  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_gray_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_sync_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.fifo_rptr_sync_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.fifo_wptr_gray_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.fifo_wptr_gray_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.fifo_wptr_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.fifo_wptr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.storage   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_tx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_tx_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.pos  == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.pos   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.rptr == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.rptr  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.sram_rdata_q == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.sram_rdata_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.sram_req == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.sram_req  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.st   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.st    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_fwmode.u_txf_ctrl.wptr_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_fwmode.u_txf_ctrl.wptr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.a_rvalid_sram_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.a_rvalid_sram_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.b_rvalid_sram_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.b_rvalid_sram_q   &&
  //      top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o   == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o    &&
 //       top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o   == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o    &&
 //       top_level_upec.top_earlgrey_1.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.mem == top_level_upec.top_earlgrey_2.u_spi_device.u_memory_2p.u_mem.gen_generic.u_impl_generic.mem  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_p2s.cnt    == top_level_upec.top_earlgrey_2.u_spi_device.u_p2s.cnt &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_p2s.io_mode    == top_level_upec.top_earlgrey_2.u_spi_device.u_p2s.io_mode &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_p2s.out_shift  == top_level_upec.top_earlgrey_2.u_spi_device.u_p2s.out_shift   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_p2s.tx_state   == top_level_upec.top_earlgrey_2.u_spi_device.u_p2s.tx_state    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.addr_phase_outclk  == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.addr_phase_outclk   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.addrcnt    == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.addrcnt &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.addrcnt_outclk == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.addrcnt_outclk  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.bitcnt == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.bitcnt  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.cmd_filter == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.cmd_filter  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.cmd_info   == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.cmd_info    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.cmd_info_7th   == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.cmd_info_7th    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.csb_deassert   == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.csb_deassert    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.csb_deassert_outclk    == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.csb_deassert_outclk &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.dummycnt   == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.dummycnt    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.host_s_en_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.host_s_en_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.mailbox_hit    == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.mailbox_hit &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.opcode == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.opcode  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.passthrough_s_en   == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.passthrough_s_en    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_passthrough.st == top_level_upec.top_earlgrey_2.u_spi_device.u_passthrough.st  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.addr_q == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.addr_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.bitcnt == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.bitcnt  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.dummycnt   == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.dummycnt    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.fifo_byteoffset    == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.fifo_byteoffset &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.main_st    == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.main_st &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.p2s_byte_o == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.p2s_byte_o  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.p2s_valid_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.p2s_valid_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.readbuf_idx    == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.readbuf_idx &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.fifo_rptr   == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.fifo_rptr    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.fifo_wptr   == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.fifo_wptr    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.storage == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.storage  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.under_rst   == top_level_upec.top_earlgrey_2.u_spi_device.u_readcmd.u_fifo.gen_normal_fifo.under_rst    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_addr_swap_data.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_addr_swap_data.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_addr_swap_data.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_addr_swap_data.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_addr_swap_mask.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_addr_swap_mask.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_addr_swap_mask.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_addr_swap_mask.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_addr_4b_en.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_addr_4b_en.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_addr_4b_en.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_addr_4b_en.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_cpha.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_cpha.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_cpha.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_cpha.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_cpol.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_cpol.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_cpol.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_cpol.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_rx_order.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_rx_order.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_rx_order.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_rx_order.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_timer_v.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_timer_v.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_timer_v.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_timer_v.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_tx_order.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_tx_order.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cfg_tx_order.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cfg_tx_order.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_0.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_0.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_0.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_0.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_1.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_1.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_1.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_1.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_10.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_10.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_10.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_10.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_11.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_11.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_11.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_11.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_12.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_12.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_12.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_12.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_13.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_13.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_13.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_13.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_14.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_14.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_14.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_14.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_15.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_15.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_15.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_15.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_16.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_16.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_16.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_16.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_17.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_17.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_17.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_17.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_18.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_18.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_18.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_18.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_19.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_19.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_19.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_19.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_2.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_2.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_2.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_2.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_20.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_20.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_20.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_20.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_21.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_21.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_21.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_21.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_22.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_22.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_22.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_22.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_23.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_23.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_23.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_23.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_24.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_24.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_24.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_24.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_25.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_25.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_25.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_25.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_26.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_26.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_26.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_26.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_27.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_27.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_27.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_27.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_28.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_28.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_28.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_28.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_29.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_29.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_29.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_29.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_3.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_3.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_3.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_3.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_30.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_30.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_30.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_30.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_31.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_31.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_31.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_31.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_4.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_4.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_4.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_4.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_5.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_5.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_5.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_5.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_6.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_6.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_6.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_6.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_7.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_7.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_7.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_7.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_8.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_8.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_8.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_8.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_9.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_9.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_0_filter_9.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_0_filter_9.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_32.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_32.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_32.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_32.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_33.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_33.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_33.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_33.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_34.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_34.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_34.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_34.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_35.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_35.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_35.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_35.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_36.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_36.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_36.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_36.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_37.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_37.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_37.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_37.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_38.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_38.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_38.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_38.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_39.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_39.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_39.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_39.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_40.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_40.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_40.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_40.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_41.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_41.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_41.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_41.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_42.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_42.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_42.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_42.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_43.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_43.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_43.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_43.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_44.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_44.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_44.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_44.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_45.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_45.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_45.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_45.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_46.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_46.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_46.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_46.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_47.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_47.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_47.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_47.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_48.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_48.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_48.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_48.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_49.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_49.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_49.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_49.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_50.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_50.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_50.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_50.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_51.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_51.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_51.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_51.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_52.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_52.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_52.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_52.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_53.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_53.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_53.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_53.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_54.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_54.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_54.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_54.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_55.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_55.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_55.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_55.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_56.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_56.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_56.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_56.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_57.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_57.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_57.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_57.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_58.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_58.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_58.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_58.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_59.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_59.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_59.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_59.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_60.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_60.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_60.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_60.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_61.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_61.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_61.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_61.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_62.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_62.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_62.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_62.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_63.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_63.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_1_filter_63.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_1_filter_63.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_64.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_64.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_64.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_64.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_65.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_65.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_65.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_65.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_66.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_66.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_66.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_66.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_67.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_67.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_67.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_67.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_68.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_68.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_68.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_68.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_69.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_69.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_69.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_69.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_70.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_70.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_70.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_70.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_71.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_71.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_71.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_71.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_72.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_72.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_72.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_72.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_73.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_73.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_73.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_73.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_74.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_74.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_74.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_74.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_75.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_75.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_75.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_75.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_76.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_76.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_76.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_76.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_77.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_77.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_77.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_77.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_78.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_78.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_78.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_78.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_79.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_79.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_79.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_79.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_80.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_80.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_80.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_80.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_81.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_81.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_81.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_81.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_82.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_82.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_82.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_82.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_83.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_83.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_83.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_83.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_84.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_84.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_84.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_84.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_85.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_85.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_85.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_85.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_86.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_86.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_86.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_86.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_87.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_87.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_87.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_87.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_88.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_88.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_88.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_88.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_89.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_89.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_89.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_89.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_90.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_90.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_90.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_90.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_91.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_91.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_91.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_91.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_92.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_92.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_92.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_92.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_93.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_93.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_93.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_93.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_94.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_94.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_94.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_94.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_95.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_95.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_2_filter_95.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_2_filter_95.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_100.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_100.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_100.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_100.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_101.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_101.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_101.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_101.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_102.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_102.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_102.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_102.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_103.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_103.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_103.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_103.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_104.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_104.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_104.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_104.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_105.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_105.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_105.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_105.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_106.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_106.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_106.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_106.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_107.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_107.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_107.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_107.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_108.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_108.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_108.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_108.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_109.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_109.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_109.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_109.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_110.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_110.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_110.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_110.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_111.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_111.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_111.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_111.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_112.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_112.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_112.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_112.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_113.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_113.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_113.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_113.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_114.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_114.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_114.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_114.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_115.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_115.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_115.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_115.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_116.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_116.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_116.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_116.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_117.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_117.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_117.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_117.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_118.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_118.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_118.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_118.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_119.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_119.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_119.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_119.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_120.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_120.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_120.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_120.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_121.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_121.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_121.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_121.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_122.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_122.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_122.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_122.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_123.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_123.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_123.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_123.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_124.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_124.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_124.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_124.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_125.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_125.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_125.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_125.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_126.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_126.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_126.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_126.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_127.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_127.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_127.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_127.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_96.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_96.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_96.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_96.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_97.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_97.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_97.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_97.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_98.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_98.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_98.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_98.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_99.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_99.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_3_filter_99.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_3_filter_99.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_128.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_128.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_128.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_128.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_129.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_129.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_129.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_129.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_130.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_130.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_130.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_130.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_131.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_131.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_131.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_131.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_132.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_132.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_132.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_132.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_133.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_133.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_133.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_133.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_134.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_134.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_134.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_134.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_135.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_135.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_135.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_135.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_136.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_136.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_136.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_136.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_137.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_137.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_137.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_137.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_138.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_138.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_138.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_138.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_139.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_139.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_139.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_139.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_140.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_140.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_140.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_140.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_141.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_141.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_141.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_141.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_142.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_142.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_142.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_142.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_143.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_143.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_143.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_143.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_144.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_144.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_144.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_144.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_145.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_145.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_145.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_145.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_146.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_146.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_146.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_146.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_147.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_147.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_147.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_147.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_148.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_148.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_148.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_148.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_149.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_149.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_149.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_149.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_150.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_150.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_150.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_150.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_151.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_151.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_151.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_151.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_152.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_152.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_152.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_152.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_153.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_153.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_153.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_153.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_154.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_154.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_154.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_154.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_155.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_155.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_155.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_155.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_156.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_156.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_156.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_156.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_157.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_157.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_157.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_157.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_158.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_158.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_158.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_158.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_159.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_159.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_4_filter_159.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_4_filter_159.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_160.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_160.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_160.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_160.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_161.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_161.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_161.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_161.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_162.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_162.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_162.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_162.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_163.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_163.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_163.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_163.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_164.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_164.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_164.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_164.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_165.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_165.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_165.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_165.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_166.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_166.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_166.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_166.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_167.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_167.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_167.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_167.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_168.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_168.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_168.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_168.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_169.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_169.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_169.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_169.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_170.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_170.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_170.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_170.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_171.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_171.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_171.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_171.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_172.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_172.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_172.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_172.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_173.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_173.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_173.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_173.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_174.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_174.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_174.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_174.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_175.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_175.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_175.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_175.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_176.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_176.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_176.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_176.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_177.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_177.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_177.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_177.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_178.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_178.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_178.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_178.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_179.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_179.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_179.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_179.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_180.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_180.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_180.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_180.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_181.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_181.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_181.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_181.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_182.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_182.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_182.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_182.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_183.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_183.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_183.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_183.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_184.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_184.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_184.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_184.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_185.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_185.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_185.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_185.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_186.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_186.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_186.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_186.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_187.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_187.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_187.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_187.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_188.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_188.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_188.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_188.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_189.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_189.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_189.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_189.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_190.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_190.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_190.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_190.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_191.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_191.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_5_filter_191.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_5_filter_191.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_192.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_192.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_192.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_192.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_193.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_193.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_193.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_193.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_194.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_194.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_194.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_194.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_195.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_195.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_195.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_195.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_196.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_196.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_196.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_196.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_197.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_197.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_197.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_197.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_198.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_198.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_198.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_198.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_199.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_199.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_199.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_199.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_200.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_200.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_200.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_200.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_201.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_201.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_201.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_201.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_202.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_202.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_202.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_202.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_203.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_203.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_203.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_203.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_204.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_204.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_204.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_204.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_205.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_205.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_205.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_205.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_206.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_206.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_206.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_206.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_207.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_207.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_207.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_207.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_208.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_208.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_208.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_208.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_209.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_209.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_209.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_209.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_210.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_210.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_210.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_210.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_211.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_211.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_211.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_211.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_212.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_212.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_212.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_212.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_213.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_213.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_213.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_213.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_214.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_214.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_214.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_214.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_215.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_215.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_215.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_215.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_216.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_216.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_216.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_216.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_217.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_217.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_217.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_217.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_218.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_218.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_218.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_218.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_219.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_219.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_219.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_219.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_220.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_220.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_220.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_220.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_221.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_221.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_221.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_221.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_222.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_222.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_222.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_222.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_223.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_223.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_6_filter_223.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_6_filter_223.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_224.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_224.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_224.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_224.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_225.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_225.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_225.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_225.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_226.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_226.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_226.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_226.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_227.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_227.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_227.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_227.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_228.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_228.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_228.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_228.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_229.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_229.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_229.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_229.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_230.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_230.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_230.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_230.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_231.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_231.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_231.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_231.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_232.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_232.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_232.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_232.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_233.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_233.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_233.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_233.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_234.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_234.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_234.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_234.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_235.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_235.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_235.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_235.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_236.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_236.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_236.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_236.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_237.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_237.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_237.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_237.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_238.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_238.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_238.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_238.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_239.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_239.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_239.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_239.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_240.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_240.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_240.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_240.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_241.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_241.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_241.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_241.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_242.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_242.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_242.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_242.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_243.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_243.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_243.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_243.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_244.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_244.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_244.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_244.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_245.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_245.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_245.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_245.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_246.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_246.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_246.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_246.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_247.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_247.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_247.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_247.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_248.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_248.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_248.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_248.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_249.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_249.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_249.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_249.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_250.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_250.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_250.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_250.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_251.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_251.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_251.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_251.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_252.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_252.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_252.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_252.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_253.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_253.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_253.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_253.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_254.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_254.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_254.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_254.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_255.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_255.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_filter_7_filter_255.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_filter_7_filter_255.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_4b_affected_0.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_4b_affected_0.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_4b_affected_0.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_4b_affected_0.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_en_0.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_en_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_en_0.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_en_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_swap_en_0.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_swap_en_0.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_addr_swap_en_0.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_addr_swap_en_0.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_dummy_en_0.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_dummy_en_0.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_dummy_en_0.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_dummy_en_0.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_dummy_size_0.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_dummy_size_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_dummy_size_0.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_dummy_size_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_opcode_0.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_opcode_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_opcode_0.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_opcode_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_payload_dir_0.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_payload_dir_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_payload_dir_0.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_payload_dir_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_payload_en_0.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_payload_en_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_0_payload_en_0.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_0_payload_en_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_4b_affected_10.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_4b_affected_10.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_4b_affected_10.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_4b_affected_10.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_en_10.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_en_10.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_en_10.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_en_10.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_swap_en_10.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_swap_en_10.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_addr_swap_en_10.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_addr_swap_en_10.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_dummy_en_10.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_dummy_en_10.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_dummy_en_10.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_dummy_en_10.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_dummy_size_10.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_dummy_size_10.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_dummy_size_10.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_dummy_size_10.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_opcode_10.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_opcode_10.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_opcode_10.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_opcode_10.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_payload_dir_10.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_payload_dir_10.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_payload_dir_10.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_payload_dir_10.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_payload_en_10.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_payload_en_10.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_10_payload_en_10.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_10_payload_en_10.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_4b_affected_11.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_4b_affected_11.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_4b_affected_11.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_4b_affected_11.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_en_11.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_en_11.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_en_11.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_en_11.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_swap_en_11.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_swap_en_11.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_addr_swap_en_11.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_addr_swap_en_11.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_dummy_en_11.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_dummy_en_11.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_dummy_en_11.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_dummy_en_11.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_dummy_size_11.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_dummy_size_11.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_dummy_size_11.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_dummy_size_11.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_opcode_11.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_opcode_11.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_opcode_11.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_opcode_11.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_payload_dir_11.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_payload_dir_11.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_payload_dir_11.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_payload_dir_11.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_payload_en_11.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_payload_en_11.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_11_payload_en_11.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_11_payload_en_11.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_4b_affected_12.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_4b_affected_12.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_4b_affected_12.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_4b_affected_12.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_en_12.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_en_12.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_en_12.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_en_12.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_swap_en_12.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_swap_en_12.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_addr_swap_en_12.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_addr_swap_en_12.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_dummy_en_12.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_dummy_en_12.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_dummy_en_12.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_dummy_en_12.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_dummy_size_12.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_dummy_size_12.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_dummy_size_12.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_dummy_size_12.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_opcode_12.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_opcode_12.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_opcode_12.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_opcode_12.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_payload_dir_12.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_payload_dir_12.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_payload_dir_12.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_payload_dir_12.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_payload_en_12.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_payload_en_12.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_12_payload_en_12.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_12_payload_en_12.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_4b_affected_13.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_4b_affected_13.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_4b_affected_13.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_4b_affected_13.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_en_13.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_en_13.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_en_13.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_en_13.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_swap_en_13.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_swap_en_13.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_addr_swap_en_13.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_addr_swap_en_13.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_dummy_en_13.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_dummy_en_13.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_dummy_en_13.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_dummy_en_13.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_dummy_size_13.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_dummy_size_13.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_dummy_size_13.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_dummy_size_13.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_opcode_13.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_opcode_13.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_opcode_13.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_opcode_13.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_payload_dir_13.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_payload_dir_13.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_payload_dir_13.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_payload_dir_13.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_payload_en_13.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_payload_en_13.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_13_payload_en_13.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_13_payload_en_13.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_4b_affected_14.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_4b_affected_14.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_4b_affected_14.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_4b_affected_14.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_en_14.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_en_14.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_en_14.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_en_14.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_swap_en_14.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_swap_en_14.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_addr_swap_en_14.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_addr_swap_en_14.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_dummy_en_14.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_dummy_en_14.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_dummy_en_14.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_dummy_en_14.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_dummy_size_14.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_dummy_size_14.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_dummy_size_14.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_dummy_size_14.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_opcode_14.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_opcode_14.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_opcode_14.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_opcode_14.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_payload_dir_14.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_payload_dir_14.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_payload_dir_14.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_payload_dir_14.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_payload_en_14.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_payload_en_14.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_14_payload_en_14.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_14_payload_en_14.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_4b_affected_15.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_4b_affected_15.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_4b_affected_15.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_4b_affected_15.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_en_15.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_en_15.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_en_15.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_en_15.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_swap_en_15.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_swap_en_15.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_addr_swap_en_15.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_addr_swap_en_15.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_dummy_en_15.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_dummy_en_15.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_dummy_en_15.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_dummy_en_15.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_dummy_size_15.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_dummy_size_15.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_dummy_size_15.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_dummy_size_15.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_opcode_15.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_opcode_15.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_opcode_15.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_opcode_15.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_payload_dir_15.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_payload_dir_15.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_payload_dir_15.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_payload_dir_15.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_payload_en_15.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_payload_en_15.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_15_payload_en_15.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_15_payload_en_15.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_4b_affected_1.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_4b_affected_1.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_4b_affected_1.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_4b_affected_1.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_en_1.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_en_1.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_en_1.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_en_1.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_swap_en_1.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_swap_en_1.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_addr_swap_en_1.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_addr_swap_en_1.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_dummy_en_1.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_dummy_en_1.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_dummy_en_1.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_dummy_en_1.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_dummy_size_1.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_dummy_size_1.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_dummy_size_1.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_dummy_size_1.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_opcode_1.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_opcode_1.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_opcode_1.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_opcode_1.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_payload_dir_1.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_payload_dir_1.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_payload_dir_1.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_payload_dir_1.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_payload_en_1.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_payload_en_1.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_1_payload_en_1.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_1_payload_en_1.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_4b_affected_2.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_4b_affected_2.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_4b_affected_2.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_4b_affected_2.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_en_2.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_en_2.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_en_2.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_en_2.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_swap_en_2.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_swap_en_2.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_addr_swap_en_2.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_addr_swap_en_2.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_dummy_en_2.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_dummy_en_2.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_dummy_en_2.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_dummy_en_2.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_dummy_size_2.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_dummy_size_2.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_dummy_size_2.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_dummy_size_2.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_opcode_2.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_opcode_2.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_opcode_2.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_opcode_2.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_payload_dir_2.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_payload_dir_2.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_payload_dir_2.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_payload_dir_2.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_payload_en_2.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_payload_en_2.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_2_payload_en_2.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_2_payload_en_2.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_4b_affected_3.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_4b_affected_3.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_4b_affected_3.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_4b_affected_3.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_en_3.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_en_3.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_en_3.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_en_3.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_swap_en_3.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_swap_en_3.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_addr_swap_en_3.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_addr_swap_en_3.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_dummy_en_3.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_dummy_en_3.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_dummy_en_3.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_dummy_en_3.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_dummy_size_3.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_dummy_size_3.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_dummy_size_3.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_dummy_size_3.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_opcode_3.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_opcode_3.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_opcode_3.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_opcode_3.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_payload_dir_3.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_payload_dir_3.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_payload_dir_3.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_payload_dir_3.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_payload_en_3.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_payload_en_3.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_3_payload_en_3.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_3_payload_en_3.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_4b_affected_4.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_4b_affected_4.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_4b_affected_4.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_4b_affected_4.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_en_4.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_en_4.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_en_4.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_en_4.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_swap_en_4.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_swap_en_4.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_addr_swap_en_4.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_addr_swap_en_4.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_dummy_en_4.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_dummy_en_4.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_dummy_en_4.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_dummy_en_4.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_dummy_size_4.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_dummy_size_4.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_dummy_size_4.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_dummy_size_4.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_opcode_4.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_opcode_4.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_opcode_4.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_opcode_4.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_payload_dir_4.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_payload_dir_4.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_payload_dir_4.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_payload_dir_4.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_payload_en_4.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_payload_en_4.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_4_payload_en_4.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_4_payload_en_4.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_4b_affected_5.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_4b_affected_5.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_4b_affected_5.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_4b_affected_5.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_en_5.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_en_5.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_en_5.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_en_5.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_swap_en_5.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_swap_en_5.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_addr_swap_en_5.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_addr_swap_en_5.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_dummy_en_5.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_dummy_en_5.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_dummy_en_5.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_dummy_en_5.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_dummy_size_5.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_dummy_size_5.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_dummy_size_5.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_dummy_size_5.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_opcode_5.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_opcode_5.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_opcode_5.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_opcode_5.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_payload_dir_5.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_payload_dir_5.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_payload_dir_5.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_payload_dir_5.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_payload_en_5.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_payload_en_5.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_5_payload_en_5.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_5_payload_en_5.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_4b_affected_6.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_4b_affected_6.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_4b_affected_6.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_4b_affected_6.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_en_6.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_en_6.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_en_6.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_en_6.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_swap_en_6.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_swap_en_6.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_addr_swap_en_6.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_addr_swap_en_6.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_dummy_en_6.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_dummy_en_6.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_dummy_en_6.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_dummy_en_6.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_dummy_size_6.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_dummy_size_6.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_dummy_size_6.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_dummy_size_6.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_opcode_6.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_opcode_6.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_opcode_6.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_opcode_6.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_payload_dir_6.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_payload_dir_6.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_payload_dir_6.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_payload_dir_6.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_payload_en_6.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_payload_en_6.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_6_payload_en_6.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_6_payload_en_6.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_4b_affected_7.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_4b_affected_7.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_4b_affected_7.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_4b_affected_7.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_en_7.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_en_7.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_en_7.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_en_7.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_swap_en_7.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_swap_en_7.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_addr_swap_en_7.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_addr_swap_en_7.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_dummy_en_7.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_dummy_en_7.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_dummy_en_7.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_dummy_en_7.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_dummy_size_7.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_dummy_size_7.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_dummy_size_7.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_dummy_size_7.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_opcode_7.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_opcode_7.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_opcode_7.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_opcode_7.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_payload_dir_7.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_payload_dir_7.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_payload_dir_7.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_payload_dir_7.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_payload_en_7.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_payload_en_7.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_7_payload_en_7.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_7_payload_en_7.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_4b_affected_8.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_4b_affected_8.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_4b_affected_8.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_4b_affected_8.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_en_8.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_en_8.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_en_8.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_en_8.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_swap_en_8.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_swap_en_8.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_addr_swap_en_8.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_addr_swap_en_8.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_dummy_en_8.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_dummy_en_8.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_dummy_en_8.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_dummy_en_8.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_dummy_size_8.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_dummy_size_8.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_dummy_size_8.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_dummy_size_8.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_opcode_8.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_opcode_8.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_opcode_8.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_opcode_8.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_payload_dir_8.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_payload_dir_8.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_payload_dir_8.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_payload_dir_8.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_payload_en_8.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_payload_en_8.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_8_payload_en_8.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_8_payload_en_8.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_4b_affected_9.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_4b_affected_9.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_4b_affected_9.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_4b_affected_9.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_en_9.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_en_9.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_en_9.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_en_9.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_swap_en_9.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_swap_en_9.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_addr_swap_en_9.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_addr_swap_en_9.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_dummy_en_9.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_dummy_en_9.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_dummy_en_9.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_dummy_en_9.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_dummy_size_9.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_dummy_size_9.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_dummy_size_9.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_dummy_size_9.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_opcode_9.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_opcode_9.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_opcode_9.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_opcode_9.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_payload_dir_9.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_payload_dir_9.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_payload_dir_9.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_payload_dir_9.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_payload_en_9.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_payload_en_9.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_cmd_info_9_payload_en_9.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_cmd_info_9_payload_en_9.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_abort.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_abort.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_abort.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_abort.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_mode.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_mode.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_mode.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_mode.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_rst_rxfifo.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_rst_rxfifo.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_rst_rxfifo.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_rst_rxfifo.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_rst_txfifo.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_rst_txfifo.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_rst_txfifo.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_rst_txfifo.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_sram_clk_en.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_sram_clk_en.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_control_sram_clk_en.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_control_sram_clk_en.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_fifo_level_rxlvl.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_fifo_level_rxlvl.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_fifo_level_rxlvl.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_fifo_level_rxlvl.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_fifo_level_txlvl.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_fifo_level_txlvl.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_fifo_level_txlvl.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_fifo_level_txlvl.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxerr.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxerr.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxerr.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxerr.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxf.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxf.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxf.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxf.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxlvl.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxlvl.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxlvl.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxlvl.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxoverflow.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxoverflow.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_rxoverflow.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_rxoverflow.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_txlvl.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_txlvl.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_txlvl.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_txlvl.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_txunderflow.q    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_txunderflow.q &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_enable_txunderflow.qe   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_enable_txunderflow.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxerr.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxerr.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxerr.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxerr.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxf.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxf.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxf.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxf.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxlvl.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxlvl.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxlvl.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxlvl.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxoverflow.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxoverflow.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_rxoverflow.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_rxoverflow.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_txlvl.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_txlvl.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_txlvl.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_txlvl.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_txunderflow.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_txunderflow.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_intr_state_txunderflow.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_intr_state_txunderflow.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_addr_base.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_addr_base.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_addr_base.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_addr_base.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_addr_limit.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_addr_limit.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_addr_limit.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_addr_limit.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_ptr_rptr.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_ptr_rptr.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_ptr_rptr.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_ptr_rptr.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_ptr_wptr.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_ptr_wptr.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_rxf_ptr_wptr.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_rxf_ptr_wptr.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.dev_select_outstanding    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.dev_select_outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.err_resp.err_opcode   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.err_resp.err_opcode    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.err_resp.err_req_pending  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.err_resp.err_req_pending   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.err_resp.err_rsp_pending  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.err_resp.err_rsp_pending   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.err_resp.err_size == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.err_resp.err_size  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.err_resp.err_source   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.err_resp.err_source    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_socket.num_req_outstanding   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_socket.num_req_outstanding    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_addr_base.q  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_addr_base.q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_addr_base.qe == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_addr_base.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_addr_limit.q == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_addr_limit.q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_addr_limit.qe    == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_addr_limit.qe &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_ptr_rptr.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_ptr_rptr.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_ptr_rptr.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_ptr_rptr.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_ptr_wptr.q   == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_ptr_wptr.q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_reg.u_txf_ptr_wptr.qe  == top_level_upec.top_earlgrey_2.u_spi_device.u_reg.u_txf_ptr_wptr.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_rxf_overflow.dst_level_q   == top_level_upec.top_earlgrey_2.u_spi_device.u_rxf_overflow.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_rxf_overflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_rxf_overflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_rxf_overflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_rxf_overflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_rxf_overflow.src_level == top_level_upec.top_earlgrey_2.u_spi_device.u_rxf_overflow.src_level  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_s2p.bitcnt == top_level_upec.top_earlgrey_2.u_spi_device.u_s2p.bitcnt  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_s2p.cnt    == top_level_upec.top_earlgrey_2.u_spi_device.u_s2p.cnt &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_s2p.data_q == top_level_upec.top_earlgrey_2.u_spi_device.u_s2p.data_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sram_clk_cg.gen_generic.u_impl_generic.en_latch    == top_level_upec.top_earlgrey_2.u_spi_device.u_sram_clk_cg.gen_generic.u_impl_generic.en_latch &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_csb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_csb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_csb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_csb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_rxf.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_rxf.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_rxf.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_rxf.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_txe.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_txe.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_sync_txe.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_device.u_sync_txe.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.intg_error_q == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.intg_error_q  &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_reqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_rspfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_spi_device.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_txf_underflow.dst_level_q  == top_level_upec.top_earlgrey_2.u_spi_device.u_txf_underflow.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_txf_underflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_device.u_txf_underflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_txf_underflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_device.u_txf_underflow.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_device.u_txf_underflow.src_level    == top_level_upec.top_earlgrey_2.u_spi_device.u_txf_underflow.src_level &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.idle_q    == top_level_upec.top_earlgrey_2.u_spi_host0.idle_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.intr_hw_error.intr_o  == top_level_upec.top_earlgrey_2.u_spi_host0.intr_hw_error.intr_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.intr_hw_spi_event.intr_o  == top_level_upec.top_earlgrey_2.u_spi_host0.intr_hw_spi_event.intr_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.ready_q   == top_level_upec.top_earlgrey_2.u_spi_host0.ready_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.rx_full_q == top_level_upec.top_earlgrey_2.u_spi_host0.rx_full_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.rx_wm_q   == top_level_upec.top_earlgrey_2.u_spi_host0.rx_wm_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.tx_empty_q    == top_level_upec.top_earlgrey_2.u_spi_host0.tx_empty_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.tx_wm_q   == top_level_upec.top_earlgrey_2.u_spi_host0.tx_wm_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.cdc_req_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.cdc_req_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.command_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.command_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_ack_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_ack_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_fsm_cs == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_fsm_cs == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_req_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_req_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host0.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_csaat.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_csaat.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_csaat.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_csaat.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_direction.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_direction.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_direction.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_direction.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_len.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_len.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_len.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_len.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_speed.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_speed.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_command_speed.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_command_speed.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_clkdiv_0.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_clkdiv_0.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_clkdiv_0.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_clkdiv_0.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_cpha_0.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_cpha_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_cpha_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_cpha_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_cpol_0.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_cpol_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_cpol_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_cpol_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csnidle_0.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csnidle_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csnidle_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csnidle_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csnlead_0.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csnlead_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csnlead_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csnlead_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csntrail_0.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csntrail_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_csntrail_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_csntrail_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_fullcyc_0.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_fullcyc_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_configopts_fullcyc_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_configopts_fullcyc_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_passthru.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_passthru.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_passthru.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_passthru.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_spien.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_spien.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_spien.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_spien.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_sw_rst.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_sw_rst.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_sw_rst.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_sw_rst.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_control_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_control_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_csid.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_csid.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_csid.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_csid.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_cmdbusy.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_cmdbusy.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_cmdbusy.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_cmdbusy.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_cmdinval.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_cmdinval.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_cmdinval.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_cmdinval.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_csidinval.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_csidinval.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_csidinval.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_csidinval.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_overflow.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_overflow.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_underflow.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_underflow.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_enable_underflow.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_enable_underflow.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_cmdbusy.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_cmdbusy.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_cmdbusy.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_cmdbusy.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_cmdinval.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_cmdinval.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_cmdinval.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_cmdinval.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_csidinval.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_csidinval.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_csidinval.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_csidinval.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_overflow.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_overflow.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_underflow.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_underflow.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_error_status_underflow.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_error_status_underflow.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_idle.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_idle.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_idle.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_idle.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_ready.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_ready.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_ready.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_ready.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_rxfull.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_rxfull.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_rxfull.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_rxfull.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_rxwm.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_rxwm.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_rxwm.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_rxwm.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_txempty.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_txempty.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_txempty.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_txempty.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_txwm.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_txwm.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_event_enable_txwm.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_event_enable_txwm.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_enable_error.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_enable_error.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_enable_error.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_enable_error.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_enable_spi_event.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_enable_spi_event.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_enable_spi_event.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_enable_spi_event.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_state_error.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_state_error.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_state_error.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_state_error.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_state_spi_event.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_state_spi_event.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_intr_state_spi_event.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_intr_state_spi_event.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.dev_select_outstanding == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.dev_select_outstanding  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.err_resp.err_opcode    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.err_resp.err_opcode &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.err_resp.err_req_pending   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.err_resp.err_req_pending    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.err_resp.err_rsp_pending   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.err_resp.err_rsp_pending    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.err_resp.err_size  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.err_resp.err_size   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.err_resp.err_source    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.err_resp.err_source &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_socket.num_req_outstanding    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_socket.num_req_outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_active.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_active.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_active.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_active.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_byteorder.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_byteorder.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_byteorder.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_byteorder.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_ready.q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_ready.q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_ready.qe   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_ready.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxempty.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxempty.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxempty.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxempty.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxfull.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxfull.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxfull.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxfull.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxqd.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxqd.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxqd.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxqd.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxstall.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxstall.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxstall.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxstall.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxwm.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxwm.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_rxwm.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_rxwm.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txempty.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txempty.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txempty.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txempty.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txfull.q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txfull.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txfull.qe  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txfull.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txqd.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txqd.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txqd.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txqd.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txstall.q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txstall.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txstall.qe == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txstall.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txwm.q == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txwm.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_reg.u_status_txwm.qe    == top_level_upec.top_earlgrey_2.u_spi_host0.u_reg.u_status_txwm.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.bit_cntr_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.bit_cntr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.bit_shifting_cpha1   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.bit_shifting_cpha1    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.byte_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.byte_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.byte_ending_cpha1    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.byte_ending_cpha1 &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.byte_starting_cpha1  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.byte_starting_cpha1   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.clk_cntr_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.clk_cntr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.clkdiv_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.clkdiv_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.cmd_rd_en_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.cmd_rd_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.cmd_speed_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.cmd_speed_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.cmd_wr_en_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.cmd_wr_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.cpha_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.cpha_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.cpol_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.cpol_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csaat_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csaat_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csb_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csb_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csid_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csid_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csnidle_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csnidle_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csnlead_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csnlead_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.csntrail_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.csntrail_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.full_cyc_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.full_cyc_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.idle_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.idle_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.lead_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.lead_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.sample_en_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.sample_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.sample_en_q2 == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.sample_en_q2  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.sck_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.sck_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.spi_host_st_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.spi_host_st_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_fsm.trail_cntr_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_fsm.trail_cntr_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_merge.last_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_merge.last_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_merge.u_packer.clr_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_merge.u_packer.clr_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_merge.u_packer.data_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_merge.u_packer.data_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_merge.u_packer.depth_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_merge.u_packer.depth_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_select.u_packer.clr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_select.u_packer.clr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_select.u_packer.data_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_select.u_packer.data_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_select.u_packer.depth_q  == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_select.u_packer.depth_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_select.u_packer.gen_unpack_mode.ptr_q    == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_select.u_packer.gen_unpack_mode.ptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_shift_reg.rx_buf_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_shift_reg.rx_buf_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_shift_reg.rx_buf_valid_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_shift_reg.rx_buf_valid_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_shift_reg.sd_i_q == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_shift_reg.sd_i_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_spi_core.u_shift_reg.sr_q   == top_level_upec.top_earlgrey_2.u_spi_host0.u_spi_core.u_shift_reg.sr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host0.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host0.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host0.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host0.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.error  == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.error   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.outstanding    == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.rdata  == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.rdata   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.reqid  == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.reqid   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.reqsz  == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.reqsz   &&
        top_level_upec.top_earlgrey_1.u_spi_host0.u_window.u_adapter.rspop  == top_level_upec.top_earlgrey_2.u_spi_host0.u_window.u_adapter.rspop   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.idle_q    == top_level_upec.top_earlgrey_2.u_spi_host1.idle_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.intr_hw_error.intr_o  == top_level_upec.top_earlgrey_2.u_spi_host1.intr_hw_error.intr_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.intr_hw_spi_event.intr_o  == top_level_upec.top_earlgrey_2.u_spi_host1.intr_hw_spi_event.intr_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.ready_q   == top_level_upec.top_earlgrey_2.u_spi_host1.ready_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.rx_full_q == top_level_upec.top_earlgrey_2.u_spi_host1.rx_full_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.rx_wm_q   == top_level_upec.top_earlgrey_2.u_spi_host1.rx_wm_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.tx_empty_q    == top_level_upec.top_earlgrey_2.u_spi_host1.tx_empty_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.tx_wm_q   == top_level_upec.top_earlgrey_2.u_spi_host1.tx_wm_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.cdc_req_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.cdc_req_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.command_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.command_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_ack_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_ack_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_fsm_cs == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.dst_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_fsm_cs == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_req_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_cmd_cdc.u_sync_reqack.u_prim_sync_reqack.src_req_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_rptr    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_rptr &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_wptr    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.fifo_wptr &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.storage  == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.storage   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.under_rst    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.gen_tx_async_plus_sync.u_tx_sync_fifo.gen_normal_fifo.under_rst &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_rx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.storage    == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_spi_host1.u_data_cdc.u_tx_async_fifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_csaat.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_csaat.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_csaat.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_csaat.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_direction.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_direction.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_direction.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_direction.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_len.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_len.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_len.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_len.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_speed.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_speed.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_command_speed.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_command_speed.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_clkdiv_0.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_clkdiv_0.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_clkdiv_0.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_clkdiv_0.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_cpha_0.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_cpha_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_cpha_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_cpha_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_cpol_0.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_cpol_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_cpol_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_cpol_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csnidle_0.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csnidle_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csnidle_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csnidle_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csnlead_0.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csnlead_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csnlead_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csnlead_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csntrail_0.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csntrail_0.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_csntrail_0.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_csntrail_0.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_fullcyc_0.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_fullcyc_0.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_configopts_fullcyc_0.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_configopts_fullcyc_0.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_passthru.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_passthru.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_passthru.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_passthru.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_spien.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_spien.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_spien.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_spien.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_sw_rst.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_sw_rst.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_sw_rst.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_sw_rst.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_control_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_control_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_csid.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_csid.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_csid.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_csid.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_cmdbusy.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_cmdbusy.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_cmdbusy.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_cmdbusy.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_cmdinval.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_cmdinval.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_cmdinval.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_cmdinval.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_csidinval.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_csidinval.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_csidinval.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_csidinval.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_overflow.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_overflow.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_underflow.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_underflow.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_enable_underflow.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_enable_underflow.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_cmdbusy.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_cmdbusy.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_cmdbusy.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_cmdbusy.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_cmdinval.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_cmdinval.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_cmdinval.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_cmdinval.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_csidinval.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_csidinval.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_csidinval.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_csidinval.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_overflow.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_overflow.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_overflow.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_overflow.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_underflow.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_underflow.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_error_status_underflow.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_error_status_underflow.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_idle.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_idle.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_idle.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_idle.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_ready.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_ready.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_ready.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_ready.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_rxfull.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_rxfull.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_rxfull.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_rxfull.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_rxwm.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_rxwm.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_rxwm.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_rxwm.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_txempty.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_txempty.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_txempty.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_txempty.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_txwm.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_txwm.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_event_enable_txwm.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_event_enable_txwm.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_enable_error.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_enable_error.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_enable_error.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_enable_error.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_enable_spi_event.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_enable_spi_event.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_enable_spi_event.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_enable_spi_event.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_state_error.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_state_error.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_state_error.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_state_error.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_state_spi_event.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_state_spi_event.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_intr_state_spi_event.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_intr_state_spi_event.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.dev_select_outstanding == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.dev_select_outstanding  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.err_resp.err_opcode    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.err_resp.err_opcode &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.err_resp.err_req_pending   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.err_resp.err_req_pending    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.err_resp.err_rsp_pending   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.err_resp.err_rsp_pending    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.err_resp.err_size  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.err_resp.err_size   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.err_resp.err_source    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.err_resp.err_source &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_socket.num_req_outstanding    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_socket.num_req_outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_active.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_active.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_active.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_active.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_byteorder.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_byteorder.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_byteorder.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_byteorder.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_ready.q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_ready.q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_ready.qe   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_ready.qe    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxempty.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxempty.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxempty.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxempty.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxfull.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxfull.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxfull.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxfull.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxqd.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxqd.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxqd.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxqd.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxstall.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxstall.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxstall.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxstall.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxwm.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxwm.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_rxwm.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_rxwm.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txempty.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txempty.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txempty.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txempty.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txfull.q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txfull.q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txfull.qe  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txfull.qe   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txqd.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txqd.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txqd.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txqd.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txstall.q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txstall.q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txstall.qe == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txstall.qe  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txwm.q == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txwm.q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_reg.u_status_txwm.qe    == top_level_upec.top_earlgrey_2.u_spi_host1.u_reg.u_status_txwm.qe &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.bit_cntr_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.bit_cntr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.bit_shifting_cpha1   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.bit_shifting_cpha1    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.byte_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.byte_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.byte_ending_cpha1    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.byte_ending_cpha1 &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.byte_starting_cpha1  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.byte_starting_cpha1   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.clk_cntr_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.clk_cntr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.clkdiv_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.clkdiv_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.cmd_rd_en_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.cmd_rd_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.cmd_speed_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.cmd_speed_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.cmd_wr_en_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.cmd_wr_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.cpha_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.cpha_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.cpol_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.cpol_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csaat_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csaat_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csb_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csb_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csid_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csid_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csnidle_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csnidle_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csnlead_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csnlead_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.csntrail_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.csntrail_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.full_cyc_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.full_cyc_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.idle_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.idle_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.lead_cntr_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.lead_cntr_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.sample_en_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.sample_en_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.sample_en_q2 == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.sample_en_q2  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.sck_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.sck_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.spi_host_st_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.spi_host_st_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_fsm.trail_cntr_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_fsm.trail_cntr_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_merge.last_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_merge.last_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_merge.u_packer.clr_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_merge.u_packer.clr_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_merge.u_packer.data_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_merge.u_packer.data_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_merge.u_packer.depth_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_merge.u_packer.depth_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_select.u_packer.clr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_select.u_packer.clr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_select.u_packer.data_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_select.u_packer.data_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_select.u_packer.depth_q  == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_select.u_packer.depth_q   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_select.u_packer.gen_unpack_mode.ptr_q    == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_select.u_packer.gen_unpack_mode.ptr_q &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_shift_reg.rx_buf_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_shift_reg.rx_buf_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_shift_reg.rx_buf_valid_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_shift_reg.rx_buf_valid_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_shift_reg.sd_i_q == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_shift_reg.sd_i_q  &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_spi_core.u_shift_reg.sr_q   == top_level_upec.top_earlgrey_2.u_spi_host1.u_spi_core.u_shift_reg.sr_q    &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host1.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host1.u_sync_en_to_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host1.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_spi_host1.u_sync_stat_from_core.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.error  == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.error   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.outstanding    == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.outstanding &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.rdata  == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.rdata   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.reqid  == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.reqid   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.reqsz  == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.reqsz   &&
        top_level_upec.top_earlgrey_1.u_spi_host1.u_window.u_adapter.rspop  == top_level_upec.top_earlgrey_2.u_spi_host1.u_window.u_adapter.rspop   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.escalated_q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.escalated_q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.alert_set_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.alert_set_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.alert_test_set_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.alert_test_set_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.ping_set_q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.ping_set_q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.state_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.state_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.level_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.level_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.level_q    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.level_q &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_prim_generic_flop.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[0].u_prim_alert_sender_parity.u_prim_generic_flop.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.alert_set_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.alert_set_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.alert_test_set_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.alert_test_set_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.ping_set_q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.ping_set_q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.state_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.state_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.level_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.level_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_no_async.diff_pq   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_no_async.diff_pq    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.level_q    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.level_q &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_prim_generic_flop.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.gen_alerts[1].u_prim_alert_sender_parity.u_prim_generic_flop.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.init_q    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.init_q &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.key_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.key_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.key_req_pending_q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.key_req_pending_q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.key_seed_valid_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.key_seed_valid_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.key_valid_q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.key_valid_q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.nonce_q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.nonce_q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.parity_error_q    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.parity_error_q &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_ctrl_regwen.q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_ctrl_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_ctrl_regwen.qe    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_ctrl_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_error_address.q   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_error_address.q    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_error_address.qe  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_error_address.qe   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_exec.q    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_exec.q &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_exec.qe   == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_exec.qe    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_exec_regwen.q == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_exec_regwen.q  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_exec_regwen.qe    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_exec_regwen.qe &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_ret_aon.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_sram_ctrl_ret_aon.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.cfg_auto_block_timer    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.cfg_auto_block_timer &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_ab_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_en.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_en.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_en.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_en.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_gray_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_sync_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_rptr_sync_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_wptr_gray_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_wptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_wptr_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.fifo_wptr_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.storage  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.storage   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_auto_block_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key0_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key1_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_sel.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_cfg_key2_o_sel.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_pwrb_in_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_pwrb_in_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_autoblock.i_pwrb_in_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_autoblock.i_pwrb_in_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.cfg_combo_timer == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.cfg_combo_timer  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.cfg_debounce_timer  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.cfg_debounce_timer   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.storage    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.storage &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[0].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.storage    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.storage &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[1].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.storage    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.storage &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[2].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.storage    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.storage &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_det[3].i_cfg_combo_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[0].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[1].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[2].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_bat_disable.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_ec_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_gsc_rst.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_out[3].i_cfg_com_intr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[0].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[1].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[2].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_ac_present.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key0.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key1.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_key2.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_com_sel[3].i_cfg_com_sel_pwrb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.bat_disable_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.bat_disable_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.cfg_ec_rst_timer   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.cfg_ec_rst_timer    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.combo_det_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.combo_det_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.ec_rst_l_int   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.ec_rst_l_int    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.ec_rst_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.ec_rst_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.gsc_rst_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.gsc_rst_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.storage == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.storage  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[0].i_combo_act.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.bat_disable_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.bat_disable_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.cfg_ec_rst_timer   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.cfg_ec_rst_timer    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.combo_det_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.combo_det_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.ec_rst_l_int   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.ec_rst_l_int    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.ec_rst_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.ec_rst_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.gsc_rst_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.gsc_rst_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.storage == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.storage  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[1].i_combo_act.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.bat_disable_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.bat_disable_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.cfg_ec_rst_timer   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.cfg_ec_rst_timer    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.combo_det_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.combo_det_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.ec_rst_l_int   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.ec_rst_l_int    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.ec_rst_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.ec_rst_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.gsc_rst_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.gsc_rst_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.storage == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.storage  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[2].i_combo_act.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.bat_disable_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.bat_disable_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.cfg_ec_rst_timer   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.cfg_ec_rst_timer    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.combo_det_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.combo_det_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.ec_rst_l_int   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.ec_rst_l_int    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.ec_rst_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.ec_rst_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.gsc_rst_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.gsc_rst_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_rptr_sync_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_gray_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.fifo_wptr_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.storage == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.storage  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.i_cfg_ec_rst_pulse.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combo_act[3].i_combo_act.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer1_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer1_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer2_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer2_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer_state_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.timer_state_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.trigger_h_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.trigger_h_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.trigger_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[0].i_combo_fsm.trigger_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer1_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer1_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer2_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer2_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer_state_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.timer_state_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.trigger_h_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.trigger_h_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.trigger_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[1].i_combo_fsm.trigger_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer1_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer1_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer2_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer2_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer_state_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.timer_state_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.trigger_h_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.trigger_h_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.trigger_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[2].i_combo_fsm.trigger_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer1_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer1_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer2_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer2_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer_state_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.timer_state_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.trigger_h_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.trigger_h_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.trigger_l_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.gen_combofsm[3].i_combo_fsm.trigger_l_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.storage    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.storage &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_cfg_debounce_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.dst_level_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.src_level == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo0_intr.src_level  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.dst_level_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.src_level == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo1_intr.src_level  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.dst_level_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.src_level == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo2_intr.src_level  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.dst_level_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.src_level == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_combo3_intr.src_level  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key0_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key0_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key0_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key0_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key1_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key1_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key1_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key1_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key2_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key2_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_key2_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_key2_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_combo.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_combo.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_intr.i_sysrst_ctrl_intr_o.intr_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_intr.i_sysrst_ctrl_intr_o.intr_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_ac_present_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_ac_present_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_ac_present_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_ac_present_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_bat_disable_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_bat_disable_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_bat_disable_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_bat_disable_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key0_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key1_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_key2_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_i_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_i_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_o_inv.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_inversion.i_cfg_pwrb_o_inv.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.ac_present_intr_h2l_det_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.ac_present_intr_h2l_det_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.ac_present_intr_l2h_det_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.ac_present_intr_l2h_det_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.cfg_key_intr_timer    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.cfg_key_intr_timer &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.ec_rst_l_intr_h2l_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.ec_rst_l_intr_h2l_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.ec_rst_l_intr_l2h_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.ec_rst_l_intr_l2h_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.dst_level_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.src_level    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_h2l.src_level &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.dst_level_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.src_level    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_present_l2h.src_level &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.timer_cnt_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.timer_cnt_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.timer_state_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.timer_state_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.trigger_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ac_presentintr_fsm.trigger_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ac_present_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_ec_rst_l_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key0_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key1_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key2_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_gray_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_sync_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_rptr_sync_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_wptr_gray_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_wptr_gray_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_wptr_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.fifo_wptr_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.storage  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.storage   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_key_intr_timer.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_h2l.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_h2l.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_l2h.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_cfg_pwrb_in_l2h.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.dst_level_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.src_level  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_h2l.src_level   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.dst_level_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.src_level  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_l_l2h.src_level   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_ec_rst_lintr_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_h2l.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_in_l2h.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key0intr_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_h2l.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_in_l2h.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key1intr_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_h2l.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.dst_level_q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.src_level   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_in_l2h.src_level    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_key2intr_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.dst_level_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.src_level  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_h2l.src_level   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_int_i.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.dst_level_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.src_level  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrb_l2h.src_level   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.timer_cnt_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.timer_cnt_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.timer_state_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.timer_state_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.trigger_q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.i_pwrbintr_fsm.trigger_q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key0_intr_h2l_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key0_intr_h2l_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key0_intr_l2h_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key0_intr_l2h_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key1_intr_h2l_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key1_intr_h2l_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key1_intr_l2h_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key1_intr_l2h_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key2_intr_h2l_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key2_intr_h2l_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.key2_intr_l2h_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.key2_intr_l2h_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.pwrb_intr_h2l_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.pwrb_intr_h2l_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_keyintr.pwrb_intr_l2h_det_q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_keyintr.pwrb_intr_l2h_det_q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ac_present_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ac_present_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ac_present_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ac_present_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_bat_disable_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_ec_rst_l_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key0_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key1_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_key2_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_in_i_pin.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_in_i_pin.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_0_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_0_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_1_allow.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_1_allow.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_ov.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_ov.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_q.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_pin_vis_ovd.i_cfg_pwrb_out_q.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.intg_err_q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.intg_err_q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_auto_block_enable.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_auto_block_enable.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_auto_block_enable.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_auto_block_enable.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_debounce_timer.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_debounce_timer.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_debounce_timer.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_debounce_ctl_debounce_timer.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_sel.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_sel.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_sel.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_sel.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_value.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_value.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_value.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key0_out_value.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_sel.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_sel.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_sel.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_sel.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_value.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_value.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_value.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key1_out_value.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_sel.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_sel.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_sel.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_sel.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_value.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_value.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_value.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_auto_block_out_ctl_key2_out_value.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_0.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_0.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_0.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_0.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_1.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_1.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_1.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_1.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_2.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_2.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_2.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_2.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_3.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_3.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_3.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_det_ctl_3.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_bat_disable_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_bat_disable_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_bat_disable_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_bat_disable_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_ec_rst_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_ec_rst_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_ec_rst_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_ec_rst_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_gsc_rst_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_gsc_rst_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_gsc_rst_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_gsc_rst_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_interrupt_0.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_interrupt_0.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_interrupt_0.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_0_interrupt_0.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_bat_disable_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_bat_disable_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_bat_disable_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_bat_disable_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_ec_rst_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_ec_rst_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_ec_rst_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_ec_rst_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_gsc_rst_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_gsc_rst_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_gsc_rst_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_gsc_rst_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_interrupt_1.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_interrupt_1.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_interrupt_1.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_1_interrupt_1.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_bat_disable_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_bat_disable_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_bat_disable_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_bat_disable_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_ec_rst_2.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_ec_rst_2.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_ec_rst_2.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_ec_rst_2.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_gsc_rst_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_gsc_rst_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_gsc_rst_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_gsc_rst_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_interrupt_2.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_interrupt_2.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_interrupt_2.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_2_interrupt_2.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_bat_disable_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_bat_disable_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_bat_disable_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_bat_disable_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_ec_rst_3.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_ec_rst_3.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_ec_rst_3.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_ec_rst_3.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_gsc_rst_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_gsc_rst_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_gsc_rst_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_gsc_rst_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_interrupt_3.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_interrupt_3.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_interrupt_3.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_out_ctl_3_interrupt_3.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_ac_present_sel_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_ac_present_sel_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_ac_present_sel_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_ac_present_sel_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key0_in_sel_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key0_in_sel_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key0_in_sel_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key0_in_sel_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key1_in_sel_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key1_in_sel_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key1_in_sel_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key1_in_sel_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key2_in_sel_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key2_in_sel_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key2_in_sel_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_key2_in_sel_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_pwrb_in_sel_0.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_pwrb_in_sel_0.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_pwrb_in_sel_0.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_0_pwrb_in_sel_0.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_ac_present_sel_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_ac_present_sel_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_ac_present_sel_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_ac_present_sel_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key0_in_sel_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key0_in_sel_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key0_in_sel_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key0_in_sel_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key1_in_sel_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key1_in_sel_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key1_in_sel_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key1_in_sel_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key2_in_sel_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key2_in_sel_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key2_in_sel_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_key2_in_sel_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_pwrb_in_sel_1.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_pwrb_in_sel_1.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_pwrb_in_sel_1.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_1_pwrb_in_sel_1.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_ac_present_sel_2.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_ac_present_sel_2.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_ac_present_sel_2.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_ac_present_sel_2.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key0_in_sel_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key0_in_sel_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key0_in_sel_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key0_in_sel_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key1_in_sel_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key1_in_sel_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key1_in_sel_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key1_in_sel_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key2_in_sel_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key2_in_sel_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key2_in_sel_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_key2_in_sel_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_pwrb_in_sel_2.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_pwrb_in_sel_2.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_pwrb_in_sel_2.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_2_pwrb_in_sel_2.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_ac_present_sel_3.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_ac_present_sel_3.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_ac_present_sel_3.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_ac_present_sel_3.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key0_in_sel_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key0_in_sel_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key0_in_sel_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key0_in_sel_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key1_in_sel_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key1_in_sel_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key1_in_sel_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key1_in_sel_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key2_in_sel_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key2_in_sel_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key2_in_sel_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_key2_in_sel_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_pwrb_in_sel_3.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_pwrb_in_sel_3.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_pwrb_in_sel_3.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_com_sel_ctl_3_pwrb_in_sel_3.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo0_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo0_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo0_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo0_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo1_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo1_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo1_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo1_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo2_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo2_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo2_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo2_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo3_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo3_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo3_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_combo_intr_status_combo3_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_ec_rst_ctl.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_ec_rst_ctl.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_ec_rst_ctl.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_ec_rst_ctl.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_intr_enable.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_intr_enable.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_intr_enable.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_intr_enable.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_intr_state.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_intr_state.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_intr_state.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_intr_state.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_h2l.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_h2l.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_h2l.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_h2l.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_l2h.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_l2h.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_l2h.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ac_present_l2h.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_h2l.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_h2l.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_h2l.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_h2l.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_l2h.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_l2h.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_l2h.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_ec_rst_l_l2h.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key0_in_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key1_in_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_key2_in_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_ctl_pwrb_in_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_debounce_ctl.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_debounce_ctl.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_debounce_ctl.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_debounce_ctl.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_h2l.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_h2l.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_h2l.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_h2l.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_l2h.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_l2h.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_l2h.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ac_present_l2h.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_ec_rst_l_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_h2l.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_h2l.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_h2l.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_h2l.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_l2h.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_l2h.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_l2h.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key0_in_l2h.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_h2l.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_h2l.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_h2l.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_h2l.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_l2h.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_l2h.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_l2h.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key1_in_l2h.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_h2l.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_h2l.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_h2l.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_h2l.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_l2h.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_l2h.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_l2h.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_key2_in_l2h.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_h2l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_h2l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_h2l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_h2l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_l2h.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_l2h.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_l2h.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_intr_status_pwrb_l2h.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_ac_present.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_ac_present.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_ac_present.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_ac_present.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_bat_disable.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_bat_disable.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_bat_disable.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_bat_disable.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_in.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_in.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_in.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_in.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_out.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_out.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_out.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key0_out.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_in.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_in.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_in.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_in.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_out.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_out.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_out.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key1_out.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_in.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_in.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_in.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_in.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_out.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_out.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_out.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_key2_out.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_in.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_in.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_in.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_in.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_out.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_out.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_out.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_key_invert_ctl_pwrb_out.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_0.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_0.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_0.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_0.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_1.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_1.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_1.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_bat_disable_1.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_ec_rst_l_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key0_out_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key1_out_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_key2_out_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_0.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_0.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_0.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_0.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_1.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_1.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_1.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_allowed_ctl_pwrb_out_1.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ac_present.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ac_present.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ac_present.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ac_present.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ec_rst_l.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ec_rst_l.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ec_rst_l.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_ec_rst_l.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key0_in.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key0_in.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key0_in.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key0_in.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key1_in.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key1_in.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key1_in.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key1_in.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key2_in.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key2_in.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key2_in.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_key2_in.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_pwrb_in.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_pwrb_in.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_pwrb_in.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_in_value_pwrb_in.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_bat_disable.q   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_bat_disable.q    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_bat_disable.qe  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_bat_disable.qe   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_ec_rst_l.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_ec_rst_l.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_ec_rst_l.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_ec_rst_l.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key0_out.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key0_out.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key0_out.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key0_out.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key1_out.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key1_out.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key1_out.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key1_out.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key2_out.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key2_out.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key2_out.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_key2_out.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_pwrb_out.q  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_pwrb_out.q   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_pwrb_out.qe == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_ctl_pwrb_out.qe  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_bat_disable.q == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_bat_disable.q  &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_bat_disable.qe    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_bat_disable.qe &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_ec_rst_l.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_ec_rst_l.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_ec_rst_l.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_ec_rst_l.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key0_out.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key0_out.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key0_out.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key0_out.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key1_out.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key1_out.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key1_out.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key1_out.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key2_out.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key2_out.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key2_out.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_key2_out.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_pwrb_out.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_pwrb_out.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_pwrb_out.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_pin_out_value_pwrb_out.qe    &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.error    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.error &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.outstanding  == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.outstanding   &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.rdata    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.rdata &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.reqid    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.reqid &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.reqsz    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.reqsz &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_reg_if.rspop    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_reg_if.rspop &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_regwen.q    == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_regwen.q &&
        top_level_upec.top_earlgrey_1.u_sysrst_ctrl_aon.u_reg.u_regwen.qe   == top_level_upec.top_earlgrey_2.u_sysrst_ctrl_aon.u_reg.u_regwen.qe    &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.intg_error_q == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.intg_error_q  &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_reqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_rspfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_tl_adapter_ram_ret_aon.u_sramreqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_uart0.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_llpbk.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_llpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_llpbk.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_llpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_nco.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_nco.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_nco.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_nco.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_nf.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_nf.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_nf.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_nf.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_parity_en.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_parity_en.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_parity_en.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_parity_en.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_parity_odd.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_parity_odd.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_parity_odd.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_parity_odd.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_rx.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_rx.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_rx.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_rx.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_rxblvl.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_rxblvl.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_rxblvl.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_rxblvl.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_slpbk.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_slpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_slpbk.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_slpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_tx.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_tx.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ctrl_tx.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ctrl_tx.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_rxilvl.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_rxilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_rxilvl.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_rxilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_rxrst.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_rxrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_rxrst.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_rxrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_txilvl.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_txilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_txilvl.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_txilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_txrst.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_txrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_fifo_ctrl_txrst.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_fifo_ctrl_txrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_break_err.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_break_err.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_break_err.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_break_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_frame_err.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_frame_err.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_frame_err.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_frame_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_overflow.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_overflow.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_parity_err.q   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_parity_err.q    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_parity_err.qe  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_parity_err.qe   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_timeout.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_timeout.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_tx_empty.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_tx_empty.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_tx_empty.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_tx_empty.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_enable_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_enable_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_break_err.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_break_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_break_err.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_break_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_frame_err.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_frame_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_frame_err.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_frame_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_parity_err.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_parity_err.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_parity_err.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_parity_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_timeout.q   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_timeout.qe  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_watermark.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_tx_empty.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_tx_watermark.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_tx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_intr_state_tx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_intr_state_tx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ovrd_txen.q   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ovrd_txen.q    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ovrd_txen.qe  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ovrd_txen.qe   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ovrd_txval.q  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ovrd_txval.q   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_ovrd_txval.qe == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_ovrd_txval.qe  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_timeout_ctrl_en.q == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_timeout_ctrl_en.q  &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_timeout_ctrl_en.qe    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_timeout_ctrl_en.qe &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_timeout_ctrl_val.q    == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_timeout_ctrl_val.q &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_timeout_ctrl_val.qe   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_timeout_ctrl_val.qe    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_wdata.q   == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_wdata.q    &&
        top_level_upec.top_earlgrey_1.u_uart0.u_reg.u_wdata.qe  == top_level_upec.top_earlgrey_2.u_uart0.u_reg.u_wdata.qe   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.allzero_cnt_q   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.allzero_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.break_st_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.break_st_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_break_err.intr_o == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_break_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_frame_err.intr_o == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_frame_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_overflow.intr_o  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_overflow.intr_o   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_parity_err.intr_o    == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_parity_err.intr_o &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_rx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_rx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_tx_empty.intr_o == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_tx_empty.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.intr_hw_tx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart0.uart_core.intr_hw_tx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.nco_sum_q   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.nco_sum_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_fifo_depth_prev_q    == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_fifo_depth_prev_q &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_sync_q1  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_sync_q1   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_sync_q2  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_sync_q2   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_timeout_count_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_timeout_count_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_val_q    == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_val_q &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.rx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart0.uart_core.rx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.tx_out_q    == top_level_upec.top_earlgrey_2.u_uart0.uart_core.tx_out_q &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.tx_uart_idle_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.tx_uart_idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.tx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart0.uart_core.tx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart0.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.idle_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.rx_valid_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.rx_valid_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_rx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_rx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_tx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_tx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_tx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_tx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_tx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_tx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_tx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_tx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart0.uart_core.uart_tx.tx_q    == top_level_upec.top_earlgrey_2.u_uart0.uart_core.uart_tx.tx_q &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_uart1.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_llpbk.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_llpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_llpbk.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_llpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_nco.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_nco.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_nco.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_nco.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_nf.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_nf.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_nf.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_nf.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_parity_en.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_parity_en.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_parity_en.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_parity_en.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_parity_odd.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_parity_odd.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_parity_odd.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_parity_odd.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_rx.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_rx.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_rx.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_rx.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_rxblvl.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_rxblvl.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_rxblvl.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_rxblvl.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_slpbk.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_slpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_slpbk.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_slpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_tx.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_tx.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ctrl_tx.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ctrl_tx.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_rxilvl.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_rxilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_rxilvl.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_rxilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_rxrst.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_rxrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_rxrst.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_rxrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_txilvl.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_txilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_txilvl.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_txilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_txrst.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_txrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_fifo_ctrl_txrst.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_fifo_ctrl_txrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_break_err.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_break_err.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_break_err.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_break_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_frame_err.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_frame_err.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_frame_err.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_frame_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_overflow.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_overflow.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_parity_err.q   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_parity_err.q    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_parity_err.qe  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_parity_err.qe   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_timeout.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_timeout.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_tx_empty.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_tx_empty.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_tx_empty.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_tx_empty.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_enable_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_enable_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_break_err.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_break_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_break_err.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_break_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_frame_err.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_frame_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_frame_err.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_frame_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_parity_err.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_parity_err.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_parity_err.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_parity_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_timeout.q   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_timeout.qe  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_watermark.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_tx_empty.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_tx_watermark.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_tx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_intr_state_tx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_intr_state_tx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ovrd_txen.q   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ovrd_txen.q    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ovrd_txen.qe  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ovrd_txen.qe   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ovrd_txval.q  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ovrd_txval.q   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_ovrd_txval.qe == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_ovrd_txval.qe  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_timeout_ctrl_en.q == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_timeout_ctrl_en.q  &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_timeout_ctrl_en.qe    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_timeout_ctrl_en.qe &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_timeout_ctrl_val.q    == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_timeout_ctrl_val.q &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_timeout_ctrl_val.qe   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_timeout_ctrl_val.qe    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_wdata.q   == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_wdata.q    &&
        top_level_upec.top_earlgrey_1.u_uart1.u_reg.u_wdata.qe  == top_level_upec.top_earlgrey_2.u_uart1.u_reg.u_wdata.qe   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.allzero_cnt_q   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.allzero_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.break_st_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.break_st_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_break_err.intr_o == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_break_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_frame_err.intr_o == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_frame_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_overflow.intr_o  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_overflow.intr_o   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_parity_err.intr_o    == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_parity_err.intr_o &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_rx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_rx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_tx_empty.intr_o == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_tx_empty.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.intr_hw_tx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart1.uart_core.intr_hw_tx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.nco_sum_q   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.nco_sum_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_fifo_depth_prev_q    == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_fifo_depth_prev_q &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_sync_q1  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_sync_q1   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_sync_q2  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_sync_q2   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_timeout_count_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_timeout_count_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_val_q    == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_val_q &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.rx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart1.uart_core.rx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.tx_out_q    == top_level_upec.top_earlgrey_2.u_uart1.uart_core.tx_out_q &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.tx_uart_idle_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.tx_uart_idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.tx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart1.uart_core.tx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart1.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.idle_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.rx_valid_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.rx_valid_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_rx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_rx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_tx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_tx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_tx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_tx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_tx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_tx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_tx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_tx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart1.uart_core.uart_tx.tx_q    == top_level_upec.top_earlgrey_2.u_uart1.uart_core.uart_tx.tx_q &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_uart2.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_llpbk.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_llpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_llpbk.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_llpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_nco.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_nco.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_nco.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_nco.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_nf.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_nf.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_nf.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_nf.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_parity_en.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_parity_en.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_parity_en.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_parity_en.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_parity_odd.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_parity_odd.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_parity_odd.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_parity_odd.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_rx.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_rx.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_rx.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_rx.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_rxblvl.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_rxblvl.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_rxblvl.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_rxblvl.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_slpbk.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_slpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_slpbk.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_slpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_tx.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_tx.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ctrl_tx.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ctrl_tx.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_rxilvl.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_rxilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_rxilvl.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_rxilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_rxrst.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_rxrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_rxrst.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_rxrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_txilvl.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_txilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_txilvl.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_txilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_txrst.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_txrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_fifo_ctrl_txrst.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_fifo_ctrl_txrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_break_err.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_break_err.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_break_err.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_break_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_frame_err.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_frame_err.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_frame_err.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_frame_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_overflow.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_overflow.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_parity_err.q   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_parity_err.q    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_parity_err.qe  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_parity_err.qe   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_timeout.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_timeout.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_tx_empty.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_tx_empty.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_tx_empty.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_tx_empty.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_enable_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_enable_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_break_err.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_break_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_break_err.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_break_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_frame_err.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_frame_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_frame_err.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_frame_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_parity_err.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_parity_err.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_parity_err.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_parity_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_timeout.q   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_timeout.qe  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_watermark.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_tx_empty.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_tx_watermark.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_tx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_intr_state_tx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_intr_state_tx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ovrd_txen.q   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ovrd_txen.q    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ovrd_txen.qe  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ovrd_txen.qe   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ovrd_txval.q  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ovrd_txval.q   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_ovrd_txval.qe == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_ovrd_txval.qe  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_timeout_ctrl_en.q == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_timeout_ctrl_en.q  &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_timeout_ctrl_en.qe    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_timeout_ctrl_en.qe &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_timeout_ctrl_val.q    == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_timeout_ctrl_val.q &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_timeout_ctrl_val.qe   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_timeout_ctrl_val.qe    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_wdata.q   == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_wdata.q    &&
        top_level_upec.top_earlgrey_1.u_uart2.u_reg.u_wdata.qe  == top_level_upec.top_earlgrey_2.u_uart2.u_reg.u_wdata.qe   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.allzero_cnt_q   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.allzero_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.break_st_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.break_st_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_break_err.intr_o == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_break_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_frame_err.intr_o == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_frame_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_overflow.intr_o  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_overflow.intr_o   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_parity_err.intr_o    == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_parity_err.intr_o &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_rx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_rx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_tx_empty.intr_o == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_tx_empty.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.intr_hw_tx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart2.uart_core.intr_hw_tx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.nco_sum_q   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.nco_sum_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_fifo_depth_prev_q    == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_fifo_depth_prev_q &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_sync_q1  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_sync_q1   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_sync_q2  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_sync_q2   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_timeout_count_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_timeout_count_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_val_q    == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_val_q &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.rx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart2.uart_core.rx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.tx_out_q    == top_level_upec.top_earlgrey_2.u_uart2.uart_core.tx_out_q &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.tx_uart_idle_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.tx_uart_idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.tx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart2.uart_core.tx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart2.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.idle_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.rx_valid_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.rx_valid_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_rx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_rx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_tx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_tx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_tx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_tx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_tx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_tx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_tx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_tx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart2.uart_core.uart_tx.tx_q    == top_level_upec.top_earlgrey_2.u_uart2.uart_core.uart_tx.tx_q &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.alert_set_q   == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.alert_set_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q  == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.alert_test_set_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.ping_set_q    == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.ping_set_q &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.state_q   == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.state_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.gen_no_async.diff_pq  &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q  == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ack.level_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq    == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.gen_no_async.diff_pq &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_decode_ping.level_q  &&
        top_level_upec.top_earlgrey_1.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o   == top_level_upec.top_earlgrey_2.u_uart3.gen_alert_tx[0].u_prim_alert_sender.u_prim_generic_flop.q_o    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.intg_err_q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.intg_err_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_llpbk.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_llpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_llpbk.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_llpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_nco.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_nco.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_nco.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_nco.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_nf.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_nf.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_nf.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_nf.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_parity_en.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_parity_en.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_parity_en.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_parity_en.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_parity_odd.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_parity_odd.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_parity_odd.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_parity_odd.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_rx.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_rx.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_rx.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_rx.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_rxblvl.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_rxblvl.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_rxblvl.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_rxblvl.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_slpbk.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_slpbk.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_slpbk.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_slpbk.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_tx.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_tx.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ctrl_tx.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ctrl_tx.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_rxilvl.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_rxilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_rxilvl.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_rxilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_rxrst.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_rxrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_rxrst.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_rxrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_txilvl.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_txilvl.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_txilvl.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_txilvl.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_txrst.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_txrst.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_fifo_ctrl_txrst.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_fifo_ctrl_txrst.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_break_err.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_break_err.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_break_err.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_break_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_frame_err.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_frame_err.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_frame_err.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_frame_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_overflow.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_overflow.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_parity_err.q   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_parity_err.q    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_parity_err.qe  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_parity_err.qe   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_timeout.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_timeout.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_timeout.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_timeout.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_rx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_rx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_tx_empty.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_tx_empty.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_tx_empty.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_tx_empty.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_tx_watermark.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_tx_watermark.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_enable_tx_watermark.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_enable_tx_watermark.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_break_err.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_break_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_break_err.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_break_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_frame_err.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_frame_err.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_frame_err.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_frame_err.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_overflow.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_overflow.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_overflow.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_overflow.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_parity_err.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_parity_err.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_parity_err.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_parity_err.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_timeout.q   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_timeout.q    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_timeout.qe  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_timeout.qe   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_watermark.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_rx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_rx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_tx_empty.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_tx_empty.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_tx_empty.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_tx_empty.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_tx_watermark.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_tx_watermark.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_intr_state_tx_watermark.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_intr_state_tx_watermark.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ovrd_txen.q   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ovrd_txen.q    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ovrd_txen.qe  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ovrd_txen.qe   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ovrd_txval.q  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ovrd_txval.q   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_ovrd_txval.qe == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_ovrd_txval.qe  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.error  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.error   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.outstanding    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.outstanding &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.rdata  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.rdata   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.reqid  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.reqid   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.reqsz  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.reqsz   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_reg_if.rspop  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_reg_if.rspop   &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_timeout_ctrl_en.q == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_timeout_ctrl_en.q  &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_timeout_ctrl_en.qe    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_timeout_ctrl_en.qe &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_timeout_ctrl_val.q    == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_timeout_ctrl_val.q &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_timeout_ctrl_val.qe   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_timeout_ctrl_val.qe    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_wdata.q   == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_wdata.q    &&
        top_level_upec.top_earlgrey_1.u_uart3.u_reg.u_wdata.qe  == top_level_upec.top_earlgrey_2.u_uart3.u_reg.u_wdata.qe   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.allzero_cnt_q   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.allzero_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.break_st_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.break_st_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_break_err.intr_o == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_break_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_frame_err.intr_o == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_frame_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_overflow.intr_o  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_overflow.intr_o   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_parity_err.intr_o    == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_parity_err.intr_o &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_timeout.intr_o   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_timeout.intr_o    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_rx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_rx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_tx_empty.intr_o == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_tx_empty.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.intr_hw_tx_watermark.intr_o == top_level_upec.top_earlgrey_2.u_uart3.uart_core.intr_hw_tx_watermark.intr_o  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.nco_sum_q   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.nco_sum_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_fifo_depth_prev_q    == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_fifo_depth_prev_q &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_sync_q1  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_sync_q1   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_sync_q2  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_sync_q2   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_timeout_count_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_timeout_count_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_val_q    == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_val_q &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.rx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart3.uart_core.rx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.sync_rx.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.tx_out_q    == top_level_upec.top_earlgrey_2.u_uart3.uart_core.tx_out_q &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.tx_uart_idle_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.tx_uart_idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.tx_watermark_prev_q == top_level_upec.top_earlgrey_2.u_uart3.uart_core.tx_watermark_prev_q  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_rxfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_rptr  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.fifo_wptr  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.storage   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.storage    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst == top_level_upec.top_earlgrey_2.u_uart3.uart_core.u_uart_txfifo.gen_normal_fifo.under_rst  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.idle_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.idle_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.rx_valid_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.rx_valid_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_rx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_rx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_tx.baud_div_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_tx.baud_div_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_tx.bit_cnt_q   == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_tx.bit_cnt_q    &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_tx.sreg_q  == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_tx.sreg_q   &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_tx.tick_baud_q == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_tx.tick_baud_q  &&
        top_level_upec.top_earlgrey_1.u_uart3.uart_core.uart_tx.tx_q    == top_level_upec.top_earlgrey_2.u_uart3.uart_core.uart_tx.tx_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.aon_tgl  == top_level_upec.top_earlgrey_2.u_usbdev.aon_tgl   &&
        top_level_upec.top_earlgrey_1.u_usbdev.cdc_sys_to_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.cdc_sys_to_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.cdc_sys_to_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.cdc_sys_to_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.cdc_usb_to_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.cdc_usb_to_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.cdc_usb_to_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.cdc_usb_to_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.event_link_reset_q   == top_level_upec.top_earlgrey_2.u_usbdev.event_link_reset_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.i_usbdev_iomux.cdc_io_to_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.i_usbdev_iomux.cdc_io_to_sys.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.i_usbdev_iomux.cdc_io_to_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.i_usbdev_iomux.cdc_io_to_sys.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.i_usbdev_iomux.cdc_io_to_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.i_usbdev_iomux.cdc_io_to_usb.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.i_usbdev_iomux.cdc_io_to_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.i_usbdev_iomux.cdc_io_to_usb.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_av_empty.intr_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_av_empty.intr_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_av_overflow.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_av_overflow.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_connected.intr_o    == top_level_upec.top_earlgrey_2.u_usbdev.intr_connected.intr_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_disconnected.intr_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_disconnected.intr_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_frame.intr_o    == top_level_upec.top_earlgrey_2.u_usbdev.intr_frame.intr_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_host_lost.intr_o    == top_level_upec.top_earlgrey_2.u_usbdev.intr_host_lost.intr_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_hw_pkt_received.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_hw_pkt_received.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_hw_pkt_sent.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_hw_pkt_sent.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_in_err.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_in_err.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_out_err.intr_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_out_err.intr_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_reset.intr_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_reset.intr_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_resume.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_resume.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_link_suspend.intr_o == top_level_upec.top_earlgrey_2.u_usbdev.intr_link_suspend.intr_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_bitstuff_err.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_bitstuff_err.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_crc_err.intr_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_crc_err.intr_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_full.intr_o  == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_full.intr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.intr_rx_pid_err.intr_o   == top_level_upec.top_earlgrey_2.u_usbdev.intr_rx_pid_err.intr_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_av_empty.dst_level_q  == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_av_empty.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_av_empty.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_av_empty.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_av_empty.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_av_empty.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_av_empty.src_level    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_av_empty.src_level &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_frame.dst_level_q == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_frame.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_frame.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_frame.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_frame.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_frame.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_frame.src_level   == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_frame.src_level    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_bitstuff_err.dst_level_q   == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_bitstuff_err.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_bitstuff_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_bitstuff_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_bitstuff_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_bitstuff_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_bitstuff_err.src_level == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_bitstuff_err.src_level  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_crc_err.dst_level_q    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_crc_err.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_crc_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_crc_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_crc_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_crc_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_crc_err.src_level  == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_crc_err.src_level   &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_full.dst_level_q   == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_full.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_full.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_full.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_full.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_full.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_full.src_level == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_full.src_level  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_pid_err.dst_level_q    == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_pid_err.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_pid_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_pid_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_pid_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_pid_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.sync_usb_event_rx_pid_err.src_level  == top_level_upec.top_earlgrey_2.u_usbdev.sync_usb_event_rx_pid_err.src_level   &&
        top_level_upec.top_earlgrey_1.u_usbdev.syncevent.d_sync_q   == top_level_upec.top_earlgrey_2.u_usbdev.syncevent.d_sync_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.syncevent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.syncevent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.syncevent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.syncevent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.tgl_sync_d1  == top_level_upec.top_earlgrey_2.u_usbdev.tgl_sync_d1   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.a_rvalid_sram_q  == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.a_rvalid_sram_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.b_rvalid_sram_q  == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.b_rvalid_sram_q   &&
  //      top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o   == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.a_rdata_o    &&
  //      top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o   == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.b_rdata_o    &&
  //      top_level_upec.top_earlgrey_1.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.mem == top_level_upec.top_earlgrey_2.u_usbdev.u_memory_2p.u_mem.gen_generic.u_impl_generic.mem  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.intg_err_q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.intg_err_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_avbuffer.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_avbuffer.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_avbuffer.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_avbuffer.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_buffer_0.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_buffer_0.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_buffer_0.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_buffer_0.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_pend_0.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_pend_0.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_pend_0.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_pend_0.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_rdy_0.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_rdy_0.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_rdy_0.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_rdy_0.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_size_0.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_size_0.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_0_size_0.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_0_size_0.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_buffer_10.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_buffer_10.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_buffer_10.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_buffer_10.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_pend_10.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_pend_10.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_pend_10.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_pend_10.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_rdy_10.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_rdy_10.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_rdy_10.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_rdy_10.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_size_10.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_size_10.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_10_size_10.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_10_size_10.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_buffer_11.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_buffer_11.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_buffer_11.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_buffer_11.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_pend_11.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_pend_11.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_pend_11.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_pend_11.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_rdy_11.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_rdy_11.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_rdy_11.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_rdy_11.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_size_11.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_size_11.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_11_size_11.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_11_size_11.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_buffer_1.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_buffer_1.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_buffer_1.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_buffer_1.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_pend_1.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_pend_1.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_pend_1.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_pend_1.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_rdy_1.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_rdy_1.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_rdy_1.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_rdy_1.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_size_1.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_size_1.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_1_size_1.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_1_size_1.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_buffer_2.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_buffer_2.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_buffer_2.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_buffer_2.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_pend_2.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_pend_2.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_pend_2.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_pend_2.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_rdy_2.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_rdy_2.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_rdy_2.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_rdy_2.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_size_2.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_size_2.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_2_size_2.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_2_size_2.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_buffer_3.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_buffer_3.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_buffer_3.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_buffer_3.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_pend_3.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_pend_3.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_pend_3.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_pend_3.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_rdy_3.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_rdy_3.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_rdy_3.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_rdy_3.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_size_3.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_size_3.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_3_size_3.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_3_size_3.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_buffer_4.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_buffer_4.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_buffer_4.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_buffer_4.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_pend_4.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_pend_4.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_pend_4.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_pend_4.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_rdy_4.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_rdy_4.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_rdy_4.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_rdy_4.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_size_4.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_size_4.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_4_size_4.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_4_size_4.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_buffer_5.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_buffer_5.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_buffer_5.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_buffer_5.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_pend_5.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_pend_5.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_pend_5.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_pend_5.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_rdy_5.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_rdy_5.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_rdy_5.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_rdy_5.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_size_5.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_size_5.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_5_size_5.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_5_size_5.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_buffer_6.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_buffer_6.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_buffer_6.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_buffer_6.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_pend_6.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_pend_6.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_pend_6.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_pend_6.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_rdy_6.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_rdy_6.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_rdy_6.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_rdy_6.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_size_6.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_size_6.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_6_size_6.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_6_size_6.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_buffer_7.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_buffer_7.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_buffer_7.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_buffer_7.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_pend_7.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_pend_7.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_pend_7.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_pend_7.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_rdy_7.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_rdy_7.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_rdy_7.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_rdy_7.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_size_7.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_size_7.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_7_size_7.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_7_size_7.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_buffer_8.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_buffer_8.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_buffer_8.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_buffer_8.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_pend_8.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_pend_8.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_pend_8.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_pend_8.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_rdy_8.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_rdy_8.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_rdy_8.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_rdy_8.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_size_8.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_size_8.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_8_size_8.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_8_size_8.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_buffer_9.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_buffer_9.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_buffer_9.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_buffer_9.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_pend_9.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_pend_9.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_pend_9.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_pend_9.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_rdy_9.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_rdy_9.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_rdy_9.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_rdy_9.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_size_9.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_size_9.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_configin_9_size_9.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_configin_9_size_9.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_0.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_0.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_0.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_0.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_1.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_1.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_1.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_1.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_10.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_10.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_10.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_10.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_11.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_11.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_11.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_11.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_2.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_2.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_2.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_2.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_3.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_3.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_3.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_3.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_4.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_4.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_4.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_4.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_5.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_5.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_5.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_5.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_6.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_6.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_6.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_6.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_7.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_7.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_7.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_7.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_8.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_8.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_8.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_8.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_9.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_9.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_data_toggle_clear_clear_9.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_data_toggle_clear_clear_9.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_0.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_0.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_0.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_0.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_1.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_1.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_1.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_1.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_10.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_10.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_10.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_10.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_11.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_11.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_11.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_11.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_2.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_2.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_2.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_2.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_3.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_3.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_3.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_3.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_4.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_4.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_4.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_4.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_5.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_5.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_5.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_5.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_6.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_6.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_6.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_6.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_7.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_7.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_7.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_7.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_8.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_8.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_8.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_8.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_9.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_9.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_in_sent_sent_9.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_in_sent_sent_9.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_av_empty.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_av_empty.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_av_empty.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_av_empty.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_av_overflow.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_av_overflow.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_av_overflow.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_av_overflow.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_connected.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_connected.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_connected.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_connected.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_disconnected.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_disconnected.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_disconnected.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_disconnected.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_frame.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_frame.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_frame.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_frame.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_host_lost.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_host_lost.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_host_lost.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_host_lost.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_in_err.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_in_err.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_in_err.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_in_err.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_out_err.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_out_err.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_out_err.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_out_err.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_reset.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_reset.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_reset.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_reset.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_resume.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_resume.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_resume.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_resume.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_suspend.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_suspend.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_link_suspend.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_link_suspend.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_pkt_received.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_pkt_received.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_pkt_received.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_pkt_received.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_pkt_sent.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_pkt_sent.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_pkt_sent.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_pkt_sent.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_bitstuff_err.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_bitstuff_err.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_bitstuff_err.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_bitstuff_err.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_crc_err.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_crc_err.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_crc_err.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_crc_err.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_full.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_full.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_full.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_full.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_pid_err.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_pid_err.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_enable_rx_pid_err.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_enable_rx_pid_err.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_av_empty.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_av_empty.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_av_empty.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_av_empty.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_av_overflow.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_av_overflow.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_av_overflow.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_av_overflow.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_connected.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_connected.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_connected.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_connected.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_disconnected.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_disconnected.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_disconnected.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_disconnected.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_frame.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_frame.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_frame.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_frame.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_host_lost.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_host_lost.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_host_lost.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_host_lost.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_in_err.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_in_err.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_in_err.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_in_err.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_out_err.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_out_err.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_out_err.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_out_err.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_reset.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_reset.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_reset.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_reset.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_resume.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_resume.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_resume.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_resume.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_suspend.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_suspend.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_link_suspend.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_link_suspend.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_pkt_received.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_pkt_received.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_pkt_received.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_pkt_received.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_pkt_sent.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_pkt_sent.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_pkt_sent.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_pkt_sent.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_bitstuff_err.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_bitstuff_err.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_bitstuff_err.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_bitstuff_err.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_crc_err.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_crc_err.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_crc_err.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_crc_err.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_full.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_full.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_full.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_full.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_pid_err.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_pid_err.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_intr_state_rx_pid_err.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_intr_state_rx_pid_err.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_0.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_0.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_0.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_0.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_1.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_1.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_1.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_1.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_10.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_10.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_10.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_10.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_11.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_11.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_11.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_11.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_2.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_2.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_2.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_2.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_3.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_3.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_3.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_3.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_4.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_4.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_4.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_4.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_5.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_5.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_5.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_5.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_6.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_6.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_6.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_6.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_7.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_7.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_7.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_7.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_8.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_8.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_8.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_8.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_9.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_9.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_iso_iso_9.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_iso_iso_9.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_eop_single_bit.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_eop_single_bit.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_eop_single_bit.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_eop_single_bit.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_override_pwr_sense_en.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_override_pwr_sense_en.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_override_pwr_sense_en.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_override_pwr_sense_en.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_override_pwr_sense_val.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_override_pwr_sense_val.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_override_pwr_sense_val.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_override_pwr_sense_val.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_pinflip.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_pinflip.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_pinflip.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_pinflip.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_rx_differential_mode.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_rx_differential_mode.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_rx_differential_mode.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_rx_differential_mode.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_tx_differential_mode.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_tx_differential_mode.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_tx_differential_mode.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_tx_differential_mode.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_tx_osc_test_mode.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_tx_osc_test_mode.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_tx_osc_test_mode.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_tx_osc_test_mode.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_usb_ref_disable.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_usb_ref_disable.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_config_usb_ref_disable.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_config_usb_ref_disable.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_d_o.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_d_o.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_d_o.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_d_o.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dn_o.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dn_o.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dn_o.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dn_o.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dn_pullup_en_o.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dn_pullup_en_o.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dn_pullup_en_o.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dn_pullup_en_o.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dp_o.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dp_o.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dp_o.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dp_o.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dp_pullup_en_o.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dp_pullup_en_o.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_dp_pullup_en_o.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_dp_pullup_en_o.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_en.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_en.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_en.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_en.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_oe_o.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_oe_o.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_oe_o.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_oe_o.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_se0_o.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_se0_o.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_se0_o.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_se0_o.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_suspend_o.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_suspend_o.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_suspend_o.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_suspend_o.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_tx_mode_se_o.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_tx_mode_se_o.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_phy_pins_drive_tx_mode_se_o.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_phy_pins_drive_tx_mode_se_o.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.error == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.error  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.outstanding   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.outstanding    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.rdata == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.rdata  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.reqid == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.reqid  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.reqsz == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.reqsz  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_reg_if.rspop == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_reg_if.rspop  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_0.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_0.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_0.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_0.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_1.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_1.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_1.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_1.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_10.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_10.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_10.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_10.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_11.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_11.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_11.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_11.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_2.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_2.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_2.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_2.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_3.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_3.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_3.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_3.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_4.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_4.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_4.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_4.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_5.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_5.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_5.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_5.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_6.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_6.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_6.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_6.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_7.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_7.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_7.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_7.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_8.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_8.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_8.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_8.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_9.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_9.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_out_out_9.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_out_out_9.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_0.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_0.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_0.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_0.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_1.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_1.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_1.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_1.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_10.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_10.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_10.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_10.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_11.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_11.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_11.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_11.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_2.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_2.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_2.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_2.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_3.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_3.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_3.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_3.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_4.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_4.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_4.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_4.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_5.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_5.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_5.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_5.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_6.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_6.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_6.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_6.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_7.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_7.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_7.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_7.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_8.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_8.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_8.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_8.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_9.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_9.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_rxenable_setup_setup_9.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_rxenable_setup_setup_9.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.dev_select_outstanding    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.dev_select_outstanding &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.err_resp.err_opcode   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.err_resp.err_opcode    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.err_resp.err_req_pending  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.err_resp.err_req_pending   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.err_resp.err_rsp_pending  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.err_resp.err_rsp_pending   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.err_resp.err_size == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.err_resp.err_size  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.err_resp.err_source   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.err_resp.err_source    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_socket.num_req_outstanding   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_socket.num_req_outstanding    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_0.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_0.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_0.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_0.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_1.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_1.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_1.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_1.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_10.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_10.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_10.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_10.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_11.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_11.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_11.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_11.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_2.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_2.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_2.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_2.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_3.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_3.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_3.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_3.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_4.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_4.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_4.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_4.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_5.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_5.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_5.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_5.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_6.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_6.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_6.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_6.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_7.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_7.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_7.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_7.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_8.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_8.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_8.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_8.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_9.q  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_9.q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_stall_stall_9.qe == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_stall_stall_9.qe  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_usbctrl_device_address.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_usbctrl_device_address.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_usbctrl_device_address.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_usbctrl_device_address.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_usbctrl_enable.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_usbctrl_enable.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_usbctrl_enable.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_usbctrl_enable.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_config_wake_ack.q   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_config_wake_ack.q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_config_wake_ack.qe  == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_config_wake_ack.qe   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_config_wake_en.q    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_config_wake_en.q &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_config_wake_en.qe   == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_config_wake_en.qe    &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_debug.q == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_debug.q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_reg.u_wake_debug.qe    == top_level_upec.top_earlgrey_2.u_usbdev.u_reg.u_wake_debug.qe &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tgl_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.u_tgl_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tgl_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.u_tgl_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.intg_error_q == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.intg_error_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_reqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_rspfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_rptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.fifo_wptr   &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.storage    == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.storage &&
        top_level_upec.top_earlgrey_1.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.under_rst  == top_level_upec.top_earlgrey_2.u_usbdev.u_tlul2sram.u_sramreqfifo.gen_normal_fifo.under_rst   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usb_out_of_rst_o == top_level_upec.top_earlgrey_2.u_usbdev.usb_out_of_rst_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usb_ref_val_q    == top_level_upec.top_earlgrey_2.u_usbdev.usb_ref_val_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.storage    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.storage &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_avfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_avfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_data_toggle_clear.dst_level_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_data_toggle_clear.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_data_toggle_clear.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_data_toggle_clear.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_data_toggle_clear.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_data_toggle_clear.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_data_toggle_clear.src_level   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_data_toggle_clear.src_level    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_devclr.dst_level_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_devclr.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_devclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_devclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_devclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_devclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_devclr.src_level  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_devclr.src_level   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.av_rready_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.av_rready_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.frame_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.frame_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.ns_cnt   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.ns_cnt    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.out_max_used_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.out_max_used_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.pkt_start_rd == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.pkt_start_rd  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.std_write_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.std_write_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.data_toggle_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.data_toggle_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.ep_impl_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.ep_impl_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_current_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_current_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_data_get_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_data_get_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_get_addr_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_get_addr_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_newpkt_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_newpkt_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_rollback_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_ep_rollback_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_xfr_state    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.in_xfr_state &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.tx_data_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_in_pe.tx_data_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.current_xfer_setup_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.current_xfer_setup_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.data_toggle_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.data_toggle_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.ep_impl_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.ep_impl_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.nak_out_transfer   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.nak_out_transfer    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_current_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_current_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_data_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_data_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_data_put_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_data_put_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_newpkt_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_newpkt_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_put_addr_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_put_addr_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_setup_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_ep_setup_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_xfr_state  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_nb_out_pe.out_xfr_state   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.addr_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.addr_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bit_phase_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bit_phase_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bitstuff_error_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bitstuff_error_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bitstuff_history_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.bitstuff_history_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.crc16_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.crc16_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.crc5_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.crc5_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.diff_state_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.diff_state_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.endp_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.endp_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.frame_num_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.frame_num_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.full_pid_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.full_pid_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_history_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_history_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_state_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_state_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_state_qq == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.line_state_qq  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.packet_valid_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.packet_valid_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.rx_data_buffer_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.rx_data_buffer_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.token_payload_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_rx.token_payload_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bit_count_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bit_count_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bit_history_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bit_history_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q2   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q2    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q3   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q3    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q4   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.bitstuff_q4    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.byte_strobe_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.byte_strobe_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.crc16_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.crc16_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.data_payload_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.data_payload_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.data_shift_reg_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.data_shift_reg_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.dp_eop_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.dp_eop_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.oe_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.oe_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.oe_shift_reg_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.oe_shift_reg_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.out_state_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.out_state_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.pid_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.pid_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.se0_shift_reg_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.se0_shift_reg_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.state_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.state_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.tx_data_get_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.tx_data_get_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.usb_d_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.usb_d_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.usb_se0_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usb_fs_nb_pe.u_usb_fs_tx.usb_se0_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_pwr_sense.stored_value_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_pwr_sense.stored_value_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_pwr_sense.stored_vector_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_pwr_sense.stored_vector_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_se0.stored_value_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_se0.stored_value_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_se0.stored_vector_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.filter_se0.stored_vector_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.host_presence_timer   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.host_presence_timer    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_inac_state_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_inac_state_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_inac_timer_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_inac_timer_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_rst_state_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_rst_state_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_rst_timer_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_rst_timer_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_state_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.u_usbdev_linkstate.link_state_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_impl.wdata    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_impl.wdata &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_outrdyclr.dst_level_q == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_outrdyclr.dst_level_q  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_outrdyclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_outrdyclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_outrdyclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_outrdyclr.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_outrdyclr.src_level   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_outrdyclr.src_level    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rdysync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rdysync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rdysync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rdysync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_resume.dst_level_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_resume.dst_level_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_resume.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_resume.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_resume.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_resume.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_resume.src_level  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_resume.src_level   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.fifo_rptr_gray_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.fifo_rptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.fifo_rptr_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.fifo_rptr_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.fifo_rptr_sync_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.fifo_rptr_sync_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.fifo_wptr_gray_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.fifo_wptr_gray_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.fifo_wptr_q    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.fifo_wptr_q &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.storage    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.storage &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_rxfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_rxfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_setsent.dst_level_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_setsent.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_setsent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_setsent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_setsent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_setsent.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_setsent.src_level == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_setsent.src_level  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_ep_cfg.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_ep_cfg.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_ep_cfg.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_ep_cfg.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_in_err.dst_level_q   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_in_err.dst_level_q    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_in_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_in_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_in_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_in_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_in_err.src_level == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_in_err.src_level  &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_out_err.dst_level_q  == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_out_err.dst_level_q   &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_out_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_out_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_out_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_out_err.prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_out_err.src_level    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_out_err.src_level &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_phy_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_2.u_usbdev.usbdev_sync_phy_config.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o &&
        top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_phy_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o    == top_level_upec.top_earlgrey_1.u_usbdev.usbdev_sync_phy_config.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o
    );
endfunction