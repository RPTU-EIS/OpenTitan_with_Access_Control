function automatic input_equivalence_sram_ctrl_main();
    input_equivalence_sram_ctrl_main = (
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.alert_rx_i           == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.alert_rx_i            &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.sram_otp_key_i       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.sram_otp_key_i        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.sram_scr_i           == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.sram_scr_i            &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.sram_scr_init_i      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.sram_scr_init_i       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.lc_escalate_en_i     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.lc_escalate_en_i      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.lc_hw_debug_en_i     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.lc_hw_debug_en_i      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.otp_en_sram_ifetch_i == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.otp_en_sram_ifetch_i  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.intg_error_i         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.intg_error_i          &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.tl_i                 == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.tl_i                  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.clk_i                == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.clk_i                 &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.clk_otp_i            == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.clk_otp_i             &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.rst_ni               == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.rst_ni                &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.rst_otp_ni           == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.rst_otp_ni
    );
endfunction

function automatic output_equivalence_sram_ctrl_main();
    output_equivalence_sram_ctrl_main = (
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.sram_otp_key_o       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.sram_otp_key_o        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.sram_scr_o           == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.sram_scr_o            &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.sram_scr_init_o      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.sram_scr_init_o       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.en_ifetch_o          == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.en_ifetch_o           &&
//        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.tl_o                 == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.tl_o                  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.alert_tx_o           == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.alert_tx_o
    );
endfunction

function automatic visible_soc_state_equivalence_sram_ctrl_main();
    visible_soc_state_equivalence_sram_ctrl_main = (
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.status_error_qs                == top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.status_error_qs                 &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.status_escalated_qs            == top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.status_escalated_qs             &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.status_scr_key_valid_qs        == top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.status_scr_key_valid_qs         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.status_scr_key_seed_valid_qs   == top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.status_scr_key_seed_valid_qs    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.exec_regwen_qs                 == top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.exec_regwen_qs                  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.exec_qs                        == top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.exec_qs                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.ctrl_regwen_qs                 == top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.ctrl_regwen_qs                  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.ctrl_renew_scr_key_qs          == top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.ctrl_renew_scr_key_qs           &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.ctrl_init_qs                   == top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.ctrl_init_qs                    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.error_address_qs               == top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.error_address_qs
    );
endfunction

function automatic micro_soc_state_equivalence_sram_ctrl_main();
    micro_soc_state_equivalence_sram_ctrl_main = (
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.escalated_q                                                                                                                                  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.escalated_q                                                                                                                                   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.alert_set_q                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.alert_set_q                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.alert_test_set_q                                                                                    == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.alert_test_set_q                                                                                     &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.ping_set_q                                                                                          == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.ping_set_q                                                                                           &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.state_q                                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.state_q                                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_nq                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_nq                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_pq                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_pq                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.state_q                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.state_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.level_q                                                                                == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.level_q                                                                                 &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_nq                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_nq                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_pq                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_pq                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.state_q                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.state_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.level_q                                                                               == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.level_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_prim_generic_flop.q_o                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_prim_generic_flop.q_o                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.alert_set_q                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.alert_set_q                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.alert_test_set_q                                                                                    == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.alert_test_set_q                                                                                     &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.ping_set_q                                                                                          == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.ping_set_q                                                                                           &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.state_q                                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.state_q                                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_nq                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_nq                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_pq                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_pq                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.state_q                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.state_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.level_q                                                                                == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.level_q                                                                                 &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_nq                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_nq                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_pq                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_pq                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.state_q                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.state_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.level_q                                                                               == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.level_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_prim_generic_flop.q_o                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_prim_generic_flop.q_o                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.init_q                                                                                                                                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.init_q                                                                                                                                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.key_q                                                                                                                                        == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.key_q                                                                                                                                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.key_req_pending_q                                                                                                                            == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.key_req_pending_q                                                                                                                             &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.key_seed_valid_q                                                                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.key_seed_valid_q                                                                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.key_valid_q                                                                                                                                  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.key_valid_q                                                                                                                                   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.nonce_q                                                                                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.nonce_q                                                                                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.parity_error_q                                                                                                                               == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.parity_error_q                                                                                                                                &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                                == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                                 &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                                == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                                 &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs                                                                                        == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs                                                                                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs                                                                                        == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs                                                                                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.intg_err_q                                                                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.intg_err_q                                                                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_ctrl_regwen.q                                                                                                                        == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_ctrl_regwen.q                                                                                                                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_ctrl_regwen.qe                                                                                                                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_ctrl_regwen.qe                                                                                                                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_error_address.q                                                                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_error_address.q                                                                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_error_address.qe                                                                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_error_address.qe                                                                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_exec.q                                                                                                                               == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_exec.q                                                                                                                                &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_exec.qe                                                                                                                              == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_exec.qe                                                                                                                               &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_exec_regwen.q                                                                                                                        == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_exec_regwen.q                                                                                                                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_exec_regwen.qe                                                                                                                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_exec_regwen.qe                                                                                                                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.error                                                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.error                                                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.outstanding                                                                                                                   == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.outstanding                                                                                                                    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.rdata                                                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.rdata                                                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.reqid                                                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.reqid                                                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.reqsz                                                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.reqsz                                                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.rspop                                                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.rspop
);
endfunction

function automatic soc_state_equivalence_sram_ctrl_main();
    soc_state_equivalence_sram_ctrl_main = (
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.escalated_q                                                                                                                                  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.escalated_q                                                                                                                                   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.alert_set_q                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.alert_set_q                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.alert_test_set_q                                                                                    == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.alert_test_set_q                                                                                     &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.ping_set_q                                                                                          == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.ping_set_q                                                                                           &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.state_q                                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.state_q                                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_nq                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_nq                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_pq                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_pq                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.state_q                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.gen_async.state_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.level_q                                                                                == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ack.level_q                                                                                 &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_nq                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_nq                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_pq                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_pq                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.state_q                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.gen_async.state_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.level_q                                                                               == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_decode_ping.level_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_prim_generic_flop.q_o                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[0].u_prim_alert_sender_parity.u_prim_generic_flop.q_o                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.alert_set_q                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.alert_set_q                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.alert_test_set_q                                                                                    == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.alert_test_set_q                                                                                     &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.ping_set_q                                                                                          == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.ping_set_q                                                                                           &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.state_q                                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.state_q                                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_nq                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_nq                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_pq                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.diff_pq                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.state_q                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.gen_async.state_q                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.level_q                                                                                == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ack.level_q                                                                                 &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_nq                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_nq                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_pq                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.diff_pq                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_n.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.i_sync_p.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o  &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.state_q                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.gen_async.state_q                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.level_q                                                                               == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_decode_ping.level_q                                                                                &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_prim_generic_flop.q_o                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.gen_alerts[1].u_prim_alert_sender_parity.u_prim_generic_flop.q_o                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.init_q                                                                                                                                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.init_q                                                                                                                                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.key_q                                                                                                                                        == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.key_q                                                                                                                                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.key_req_pending_q                                                                                                                            == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.key_req_pending_q                                                                                                                             &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.key_seed_valid_q                                                                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.key_seed_valid_q                                                                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.key_valid_q                                                                                                                                  == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.key_valid_q                                                                                                                                   &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.nonce_q                                                                                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.nonce_q                                                                                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.parity_error_q                                                                                                                               == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.parity_error_q                                                                                                                                &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                                == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                                 &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                                == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_lc_sync.gen_flops.u_prim_flop_2sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                                 &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.ack_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_ack_q                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs                                                                                        == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.dst_fsm_cs                                                                                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.req_sync.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs                                                                                        == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.src_fsm_cs                                                                                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_prim_sync_reqack_data.u_prim_sync_reqack.src_req_q                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.intg_err_q                                                                                                                             == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.intg_err_q                                                                                                                              &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_ctrl_regwen.q                                                                                                                        == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_ctrl_regwen.q                                                                                                                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_ctrl_regwen.qe                                                                                                                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_ctrl_regwen.qe                                                                                                                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_error_address.q                                                                                                                      == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_error_address.q                                                                                                                       &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_error_address.qe                                                                                                                     == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_error_address.qe                                                                                                                      &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_exec.q                                                                                                                               == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_exec.q                                                                                                                                &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_exec.qe                                                                                                                              == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_exec.qe                                                                                                                               &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_exec_regwen.q                                                                                                                        == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_exec_regwen.q                                                                                                                         &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_exec_regwen.qe                                                                                                                       == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_exec_regwen.qe                                                                                                                        &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.error                                                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.error                                                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.outstanding                                                                                                                   == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.outstanding                                                                                                                    &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.rdata                                                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.rdata                                                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.reqid                                                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.reqid                                                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.reqsz                                                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.reqsz                                                                                                                          &&
        top_level_upec.top_earlgrey_1.u_sram_ctrl_main.u_reg.u_reg_if.rspop                                                                                                                         == top_level_upec.top_earlgrey_2.u_sram_ctrl_main.u_reg.u_reg_if.rspop
);
endfunction