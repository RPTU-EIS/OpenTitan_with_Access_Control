function automatic no_outstanding_reqs_to_untrusted_device_xbar_main();
    no_outstanding_reqs_to_untrusted_device_xbar_main = (
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.dev_select_outstanding           != 6'h14        &&
        top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.dev_select_outstanding           != 6'h14        &&
        !((top_level_upec.top_earlgrey_1.u_xbar_main.tl_cored_i.a_address  & 32'hfffff000)  == 32'h40300000 &&
          top_level_upec.top_earlgrey_1.u_xbar_main.tl_cored_i.a_valid)                                     &&
        !((top_level_upec.top_earlgrey_2.u_xbar_main.tl_cored_i.a_address  & 32'hfffff000)  == 32'h40300000 &&
          top_level_upec.top_earlgrey_2.u_xbar_main.tl_cored_i.a_valid)
    );
endfunction

function automatic security_enabled_xbar_main();
    security_enabled_xbar_main = (
        top_level_upec.top_earlgrey_1.u_xbar_main.master_bits_i == 1'b0 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.slave_bits_i  == 19'h7fffe
    );
endfunction

function automatic input_equivalence_xbar_main();
    input_equivalence_xbar_main = (
        top_level_upec.top_earlgrey_1.u_xbar_main.clk_main_i            == top_level_upec.top_earlgrey_2.u_xbar_main.clk_main_i             &&
        top_level_upec.top_earlgrey_1.u_xbar_main.clk_fixed_i           == top_level_upec.top_earlgrey_2.u_xbar_main.clk_fixed_i            &&
        top_level_upec.top_earlgrey_1.u_xbar_main.rst_main_ni           == top_level_upec.top_earlgrey_2.u_xbar_main.rst_main_ni            &&
        top_level_upec.top_earlgrey_1.u_xbar_main.rst_fixed_ni          == top_level_upec.top_earlgrey_2.u_xbar_main.rst_fixed_ni           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.master_bits_i         == top_level_upec.top_earlgrey_2.u_xbar_main.master_bits_i          &&
        top_level_upec.top_earlgrey_1.u_xbar_main.slave_bits_i          == top_level_upec.top_earlgrey_2.u_xbar_main.slave_bits_i           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_corei_i            == top_level_upec.top_earlgrey_2.u_xbar_main.tl_corei_i             &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_cored_i            == top_level_upec.top_earlgrey_2.u_xbar_main.tl_cored_i             &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_dm_sba_i           == top_level_upec.top_earlgrey_2.u_xbar_main.tl_dm_sba_i            &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_rom_ctrl__rom_i    == top_level_upec.top_earlgrey_2.u_xbar_main.tl_rom_ctrl__rom_i     &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_rom_ctrl__regs_i   == top_level_upec.top_earlgrey_2.u_xbar_main.tl_rom_ctrl__regs_i    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_debug_mem_i        == top_level_upec.top_earlgrey_2.u_xbar_main.tl_debug_mem_i         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_ram_main_i         == top_level_upec.top_earlgrey_2.u_xbar_main.tl_ram_main_i          &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_eflash_i           == top_level_upec.top_earlgrey_2.u_xbar_main.tl_eflash_i            &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_peri_i             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_peri_i              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_flash_ctrl__core_i == top_level_upec.top_earlgrey_2.u_xbar_main.tl_flash_ctrl__core_i  &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_flash_ctrl__prim_i == top_level_upec.top_earlgrey_2.u_xbar_main.tl_flash_ctrl__prim_i  &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_hmac_i             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_hmac_i              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_kmac_i             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_kmac_i              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_aes_i              == top_level_upec.top_earlgrey_2.u_xbar_main.tl_aes_i               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_entropy_src_i      == top_level_upec.top_earlgrey_2.u_xbar_main.tl_entropy_src_i       &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_csrng_i            == top_level_upec.top_earlgrey_2.u_xbar_main.tl_csrng_i             &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_edn0_i             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_edn0_i              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_edn1_i             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_edn1_i              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_rv_plic_i          == top_level_upec.top_earlgrey_2.u_xbar_main.tl_rv_plic_i           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_otbn_i             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_otbn_i              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_keymgr_i           == top_level_upec.top_earlgrey_2.u_xbar_main.tl_keymgr_i            &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_sram_ctrl_main_i   == top_level_upec.top_earlgrey_2.u_xbar_main.tl_sram_ctrl_main_i    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_bus_ctrl_i         == top_level_upec.top_earlgrey_2.u_xbar_main.tl_bus_ctrl_i
        );
endfunction

function automatic output_equivalence_xbar_main();
    output_equivalence_xbar_main = (
        top_level_upec.top_earlgrey_1.u_xbar_main.master_bit_peri_o     == top_level_upec.top_earlgrey_2.u_xbar_main.master_bit_peri_o       &&
        top_level_upec.top_earlgrey_1.u_xbar_main.master_bit_peri_en_o  == top_level_upec.top_earlgrey_2.u_xbar_main.master_bit_peri_en_o    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_corei_o            == top_level_upec.top_earlgrey_2.u_xbar_main.tl_corei_o              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_cored_o            == top_level_upec.top_earlgrey_2.u_xbar_main.tl_cored_o              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_dm_sba_o           == top_level_upec.top_earlgrey_2.u_xbar_main.tl_dm_sba_o             &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_rom_ctrl__rom_o    == top_level_upec.top_earlgrey_2.u_xbar_main.tl_rom_ctrl__rom_o      &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_rom_ctrl__regs_o   == top_level_upec.top_earlgrey_2.u_xbar_main.tl_rom_ctrl__regs_o     &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_debug_mem_o        == top_level_upec.top_earlgrey_2.u_xbar_main.tl_debug_mem_o          &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_ram_main_o         == top_level_upec.top_earlgrey_2.u_xbar_main.tl_ram_main_o           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_eflash_o           == top_level_upec.top_earlgrey_2.u_xbar_main.tl_eflash_o             &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_peri_o             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_peri_o               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_flash_ctrl__core_o == top_level_upec.top_earlgrey_2.u_xbar_main.tl_flash_ctrl__core_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_flash_ctrl__prim_o == top_level_upec.top_earlgrey_2.u_xbar_main.tl_flash_ctrl__prim_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_hmac_o             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_hmac_o               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_kmac_o             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_kmac_o               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_aes_o              == top_level_upec.top_earlgrey_2.u_xbar_main.tl_aes_o                &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_entropy_src_o      == top_level_upec.top_earlgrey_2.u_xbar_main.tl_entropy_src_o        &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_csrng_o            == top_level_upec.top_earlgrey_2.u_xbar_main.tl_csrng_o              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_edn0_o             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_edn0_o               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_edn1_o             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_edn1_o               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_rv_plic_o          == top_level_upec.top_earlgrey_2.u_xbar_main.tl_rv_plic_o            &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_otbn_o             == top_level_upec.top_earlgrey_2.u_xbar_main.tl_otbn_o               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_keymgr_o           == top_level_upec.top_earlgrey_2.u_xbar_main.tl_keymgr_o             &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_sram_ctrl_main_o   == top_level_upec.top_earlgrey_2.u_xbar_main.tl_sram_ctrl_main_o     &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_bus_ctrl_o         == top_level_upec.top_earlgrey_2.u_xbar_main.tl_bus_ctrl_o
    );
endfunction

function automatic core_output_equivalence_xbar_main();
    core_output_equivalence_xbar_main = (
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_corei_o    == top_level_upec.top_earlgrey_2.u_xbar_main.tl_corei_o  &&
        top_level_upec.top_earlgrey_1.u_xbar_main.tl_cored_o    == top_level_upec.top_earlgrey_2.u_xbar_main.tl_cored_o
    );
endfunction

function automatic micro_soc_state_equivalence_xbar_main();
    micro_soc_state_equivalence_xbar_main = (
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_gray_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_gray_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_q                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_sync_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_sync_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.fifo_wptr_gray_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.fifo_wptr_gray_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.fifo_wptr_q                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.fifo_wptr_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.storage                                                                      == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.storage                                                                        &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_gray_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_gray_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_q                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_sync_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_sync_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.fifo_wptr_gray_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.fifo_wptr_gray_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.fifo_wptr_q                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.fifo_wptr_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.storage                                                                      == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.storage                                                                        &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.dev_select_outstanding                                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.dev_select_outstanding                                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.err_resp.err_opcode                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.err_resp.err_opcode                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.err_resp.err_req_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.err_resp.err_req_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.err_resp.err_rsp_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.err_resp.err_rsp_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.err_resp.err_size                                                                    == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.err_resp.err_size                                                                      &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.err_resp.err_source                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.err_resp.err_source                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.num_req_outstanding                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.num_req_outstanding                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.dev_select_outstanding                                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.dev_select_outstanding                                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.err_resp.err_opcode                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.err_resp.err_opcode                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.err_resp.err_req_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.err_resp.err_req_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.err_resp.err_rsp_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.err_resp.err_rsp_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.err_resp.err_size                                                                    == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.err_resp.err_size                                                                      &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.err_resp.err_source                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.err_resp.err_source                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.num_req_outstanding                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.num_req_outstanding                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.dev_select_outstanding                                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.dev_select_outstanding                                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.err_resp.err_opcode                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.err_resp.err_opcode                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.err_resp.err_req_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.err_resp.err_req_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.err_resp.err_rsp_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.err_resp.err_rsp_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.err_resp.err_size                                                                    == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.err_resp.err_size                                                                      &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.err_resp.err_source                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.err_resp.err_source                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.fifo_rptr                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.fifo_rptr                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.fifo_wptr                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.fifo_wptr                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.storage                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.storage                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.under_rst                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.under_rst                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.fifo_rptr                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.fifo_rptr                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.fifo_wptr                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.fifo_wptr                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.storage                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.storage                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.under_rst                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.under_rst                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.num_req_outstanding                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.num_req_outstanding                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.dev_select_outstanding                                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.dev_select_outstanding                                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.err_resp.err_opcode                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.err_resp.err_opcode                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.err_resp.err_req_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.err_resp.err_req_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.err_resp.err_rsp_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.err_resp.err_rsp_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.err_resp.err_size                                                                    == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.err_resp.err_size                                                                      &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.err_resp.err_source                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.err_resp.err_source                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.num_req_outstanding                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.num_req_outstanding                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_26.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_26.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_28.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_28.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_29.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_29.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_31.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_31.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_33.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_33.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_46.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_46.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_47.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_47.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_48.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_48.gen_arb_ppc.u_reqarb.gen_normal_case.mask
    );
endfunction

function automatic soc_state_equivalence_xbar_main();
    soc_state_equivalence_xbar_main = (
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_gray_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_gray_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_q                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_sync_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.fifo_rptr_sync_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.fifo_wptr_gray_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.fifo_wptr_gray_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.fifo_wptr_q                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.fifo_wptr_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.storage                                                                      == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.storage                                                                        &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.reqfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_gray_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_gray_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_q                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_sync_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.fifo_rptr_sync_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.fifo_wptr_gray_q                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.fifo_wptr_gray_q                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.fifo_wptr_q                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.fifo_wptr_q                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.storage                                                                      == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.storage                                                                        &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.sync_rptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_1.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_asf_32.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o == top_level_upec.top_earlgrey_2.u_xbar_main.u_asf_32.rspfifo.sync_wptr.gen_generic.u_impl_generic.u_sync_2.gen_generic.u_impl_generic.q_o   &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.dev_select_outstanding                                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.dev_select_outstanding                                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.err_resp.err_opcode                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.err_resp.err_opcode                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.err_resp.err_req_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.err_resp.err_req_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.err_resp.err_rsp_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.err_resp.err_rsp_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.err_resp.err_size                                                                    == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.err_resp.err_size                                                                      &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.err_resp.err_source                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.err_resp.err_source                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_25.num_req_outstanding                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_25.num_req_outstanding                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.dev_select_outstanding                                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.dev_select_outstanding                                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.err_resp.err_opcode                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.err_resp.err_opcode                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.err_resp.err_req_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.err_resp.err_req_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.err_resp.err_rsp_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.err_resp.err_rsp_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.err_resp.err_size                                                                    == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.err_resp.err_size                                                                      &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.err_resp.err_source                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.err_resp.err_source                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_30.num_req_outstanding                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_30.num_req_outstanding                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.dev_select_outstanding                                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.dev_select_outstanding                                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.err_resp.err_opcode                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.err_resp.err_opcode                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.err_resp.err_req_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.err_resp.err_req_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.err_resp.err_rsp_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.err_resp.err_rsp_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.err_resp.err_size                                                                    == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.err_resp.err_size                                                                      &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.err_resp.err_source                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.err_resp.err_source                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.fifo_rptr                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.fifo_rptr                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.fifo_wptr                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.fifo_wptr                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.storage                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.storage                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.under_rst                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.reqfifo.gen_normal_fifo.under_rst                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.fifo_rptr                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.fifo_rptr                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.fifo_wptr                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.fifo_wptr                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.storage                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.storage                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.under_rst                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.fifo_h.rspfifo.gen_normal_fifo.under_rst                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_49.num_req_outstanding                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_49.num_req_outstanding                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.dev_select_outstanding                                                               == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.dev_select_outstanding                                                                 &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.err_resp.err_opcode                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.err_resp.err_opcode                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.err_resp.err_req_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.err_resp.err_req_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.err_resp.err_rsp_pending                                                             == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.err_resp.err_rsp_pending                                                               &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.err_resp.err_size                                                                    == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.err_resp.err_size                                                                      &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.err_resp.err_source                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.err_resp.err_source                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_s1n_50.num_req_outstanding                                                                  == top_level_upec.top_earlgrey_2.u_xbar_main.u_s1n_50.num_req_outstanding                                                                    &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_26.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_26.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_27.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_28.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_28.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_29.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_29.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_31.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_31.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_33.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_33.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_34.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_35.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_36.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_37.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_38.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_39.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_40.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_41.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_42.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_43.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_44.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.reqfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.fifo_rptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.fifo_wptr                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.storage                                         == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.storage                                           &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                       == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_45.u_devicefifo.rspfifo.gen_normal_fifo.under_rst                                         &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_46.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_46.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_47.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_47.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                              &&
        top_level_upec.top_earlgrey_1.u_xbar_main.u_sm1_48.gen_arb_ppc.u_reqarb.gen_normal_case.mask                                            == top_level_upec.top_earlgrey_2.u_xbar_main.u_sm1_48.gen_arb_ppc.u_reqarb.gen_normal_case.mask
    );
endfunction